magic
tech sky130A
magscale 1 2
timestamp 1630053115
<< checkpaint >>
rect -3932 -3932 18094 20238
<< locali >>
rect 5733 11135 5767 11305
rect 8677 10047 8711 10149
rect 8769 9911 8803 10149
rect 8711 9877 8803 9911
rect 11529 5015 11563 5185
rect 3801 2431 3835 2533
<< viali >>
rect 6745 13413 6779 13447
rect 7481 13413 7515 13447
rect 1777 13345 1811 13379
rect 10977 13345 11011 13379
rect 12173 13345 12207 13379
rect 2513 13277 2547 13311
rect 3801 13277 3835 13311
rect 4537 13277 4571 13311
rect 5181 13277 5215 13311
rect 7665 13277 7699 13311
rect 8401 13277 8435 13311
rect 9321 13277 9355 13311
rect 9505 13277 9539 13311
rect 10701 13277 10735 13311
rect 11713 13277 11747 13311
rect 11897 13277 11931 13311
rect 1961 13209 1995 13243
rect 6965 13209 6999 13243
rect 9689 13209 9723 13243
rect 11805 13209 11839 13243
rect 12035 13209 12069 13243
rect 2697 13141 2731 13175
rect 3985 13141 4019 13175
rect 4721 13141 4755 13175
rect 5365 13141 5399 13175
rect 8217 13141 8251 13175
rect 11529 13141 11563 13175
rect 11713 12937 11747 12971
rect 1777 12869 1811 12903
rect 1961 12869 1995 12903
rect 3985 12869 4019 12903
rect 10885 12869 10919 12903
rect 3433 12801 3467 12835
rect 4260 12801 4294 12835
rect 7205 12801 7239 12835
rect 7665 12801 7699 12835
rect 9045 12801 9079 12835
rect 9321 12801 9355 12835
rect 9413 12801 9447 12835
rect 11710 12801 11744 12835
rect 3893 12733 3927 12767
rect 4445 12733 4479 12767
rect 6929 12733 6963 12767
rect 7113 12733 7147 12767
rect 12173 12733 12207 12767
rect 3341 12665 3375 12699
rect 7573 12665 7607 12699
rect 9137 12665 9171 12699
rect 10609 12665 10643 12699
rect 11529 12665 11563 12699
rect 4169 12597 4203 12631
rect 9597 12597 9631 12631
rect 12081 12597 12115 12631
rect 10885 12393 10919 12427
rect 4077 12325 4111 12359
rect 11989 12257 12023 12291
rect 12265 12257 12299 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4353 12189 4387 12223
rect 9873 12189 9907 12223
rect 10793 12121 10827 12155
rect 2421 12053 2455 12087
rect 4261 12053 4295 12087
rect 9689 12053 9723 12087
rect 3249 11849 3283 11883
rect 12265 11849 12299 11883
rect 2973 11713 3007 11747
rect 3341 11713 3375 11747
rect 6544 11713 6578 11747
rect 6683 11713 6717 11747
rect 6929 11713 6963 11747
rect 10333 11713 10367 11747
rect 10793 11713 10827 11747
rect 11713 11713 11747 11747
rect 11989 11713 12023 11747
rect 12081 11713 12115 11747
rect 1409 11645 1443 11679
rect 1685 11645 1719 11679
rect 2789 11645 2823 11679
rect 11805 11645 11839 11679
rect 3065 11577 3099 11611
rect 10885 11577 10919 11611
rect 6377 11509 6411 11543
rect 6837 11509 6871 11543
rect 10149 11509 10183 11543
rect 4721 11305 4755 11339
rect 5733 11305 5767 11339
rect 12081 11305 12115 11339
rect 11345 11237 11379 11271
rect 5917 11169 5951 11203
rect 11621 11169 11655 11203
rect 4813 11101 4847 11135
rect 5733 11101 5767 11135
rect 5825 11101 5859 11135
rect 6101 11101 6135 11135
rect 6193 11101 6227 11135
rect 11069 11101 11103 11135
rect 11437 11101 11471 11135
rect 12265 11101 12299 11135
rect 6377 11033 6411 11067
rect 11161 11033 11195 11067
rect 4261 10761 4295 10795
rect 5089 10693 5123 10727
rect 5181 10693 5215 10727
rect 3985 10625 4019 10659
rect 4997 10625 5031 10659
rect 5365 10625 5399 10659
rect 3801 10557 3835 10591
rect 4353 10557 4387 10591
rect 4077 10489 4111 10523
rect 4813 10421 4847 10455
rect 2605 10217 2639 10251
rect 10057 10217 10091 10251
rect 12081 10217 12115 10251
rect 8677 10149 8711 10183
rect 2697 10013 2731 10047
rect 4537 10013 4571 10047
rect 8677 10013 8711 10047
rect 8769 10149 8803 10183
rect 1869 9945 1903 9979
rect 8953 10013 8987 10047
rect 9229 10013 9263 10047
rect 9321 10013 9355 10047
rect 9965 10013 9999 10047
rect 10977 10013 11011 10047
rect 12265 10013 12299 10047
rect 9137 9945 9171 9979
rect 1961 9877 1995 9911
rect 4445 9877 4479 9911
rect 8677 9877 8711 9911
rect 9505 9877 9539 9911
rect 11069 9877 11103 9911
rect 6653 9537 6687 9571
rect 8309 9537 8343 9571
rect 9321 9537 9355 9571
rect 8585 9469 8619 9503
rect 9045 9469 9079 9503
rect 10057 9401 10091 9435
rect 6745 9333 6779 9367
rect 7573 9333 7607 9367
rect 2881 9129 2915 9163
rect 5089 9129 5123 9163
rect 9781 9129 9815 9163
rect 1869 8993 1903 9027
rect 6009 8993 6043 9027
rect 2145 8925 2179 8959
rect 4077 8925 4111 8959
rect 4353 8925 4387 8959
rect 5733 8925 5767 8959
rect 5825 8925 5859 8959
rect 6101 8925 6135 8959
rect 9965 8925 9999 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 10057 8857 10091 8891
rect 5549 8789 5583 8823
rect 9781 8517 9815 8551
rect 8677 8449 8711 8483
rect 9597 8449 9631 8483
rect 9689 8449 9723 8483
rect 9965 8449 9999 8483
rect 8953 8381 8987 8415
rect 7941 8313 7975 8347
rect 9413 8313 9447 8347
rect 2145 7905 2179 7939
rect 2697 7905 2731 7939
rect 11989 7905 12023 7939
rect 1593 7837 1627 7871
rect 2329 7837 2363 7871
rect 12265 7837 12299 7871
rect 2605 7769 2639 7803
rect 1501 7701 1535 7735
rect 2513 7701 2547 7735
rect 1501 7497 1535 7531
rect 7481 7429 7515 7463
rect 1593 7361 1627 7395
rect 2237 7361 2271 7395
rect 3157 7361 3191 7395
rect 7757 7361 7791 7395
rect 8585 7361 8619 7395
rect 2881 7293 2915 7327
rect 7389 7293 7423 7327
rect 7941 7293 7975 7327
rect 7665 7225 7699 7259
rect 2145 7157 2179 7191
rect 3893 7157 3927 7191
rect 8493 7157 8527 7191
rect 6193 6885 6227 6919
rect 2237 6749 2271 6783
rect 2513 6749 2547 6783
rect 6377 6749 6411 6783
rect 6469 6749 6503 6783
rect 6745 6749 6779 6783
rect 7205 6749 7239 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 6561 6681 6595 6715
rect 7481 6681 7515 6715
rect 12081 6681 12115 6715
rect 1501 6613 1535 6647
rect 7757 6613 7791 6647
rect 12173 6613 12207 6647
rect 1593 6409 1627 6443
rect 2605 6409 2639 6443
rect 4537 6409 4571 6443
rect 11529 6409 11563 6443
rect 11713 6409 11747 6443
rect 7481 6341 7515 6375
rect 1409 6273 1443 6307
rect 2789 6273 2823 6307
rect 2881 6273 2915 6307
rect 3157 6273 3191 6307
rect 4534 6273 4568 6307
rect 4997 6273 5031 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 9229 6273 9263 6307
rect 10425 6273 10459 6307
rect 11710 6273 11744 6307
rect 12081 6273 12115 6307
rect 10701 6205 10735 6239
rect 12173 6205 12207 6239
rect 3065 6137 3099 6171
rect 9137 6137 9171 6171
rect 4353 6069 4387 6103
rect 4905 6069 4939 6103
rect 7205 6069 7239 6103
rect 9689 6069 9723 6103
rect 4997 5797 5031 5831
rect 4537 5729 4571 5763
rect 6469 5729 6503 5763
rect 4445 5661 4479 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 6193 5661 6227 5695
rect 7113 5661 7147 5695
rect 7205 5661 7239 5695
rect 7461 5661 7495 5695
rect 10609 5661 10643 5695
rect 10885 5661 10919 5695
rect 12173 5661 12207 5695
rect 7297 5593 7331 5627
rect 11805 5593 11839 5627
rect 11989 5593 12023 5627
rect 5457 5525 5491 5559
rect 6929 5525 6963 5559
rect 9873 5525 9907 5559
rect 3249 5321 3283 5355
rect 12265 5321 12299 5355
rect 5181 5253 5215 5287
rect 11897 5253 11931 5287
rect 3433 5185 3467 5219
rect 3525 5185 3559 5219
rect 3801 5185 3835 5219
rect 5273 5185 5307 5219
rect 6561 5185 6595 5219
rect 11529 5185 11563 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 12081 5185 12115 5219
rect 3709 5117 3743 5151
rect 6469 5049 6503 5083
rect 11529 4981 11563 5015
rect 2053 4777 2087 4811
rect 4997 4777 5031 4811
rect 9413 4777 9447 4811
rect 2605 4709 2639 4743
rect 11253 4709 11287 4743
rect 2697 4641 2731 4675
rect 2234 4573 2268 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 4073 4573 4107 4607
rect 4169 4573 4203 4607
rect 5733 4573 5767 4607
rect 6009 4573 6043 4607
rect 9505 4573 9539 4607
rect 11437 4573 11471 4607
rect 11621 4573 11655 4607
rect 11805 4573 11839 4607
rect 11529 4505 11563 4539
rect 2237 4437 2271 4471
rect 4353 4437 4387 4471
rect 3985 4233 4019 4267
rect 8953 4233 8987 4267
rect 1961 4165 1995 4199
rect 11713 4165 11747 4199
rect 11897 4165 11931 4199
rect 4077 4097 4111 4131
rect 8956 4097 8990 4131
rect 10149 4097 10183 4131
rect 10977 4097 11011 4131
rect 8493 4029 8527 4063
rect 10609 4029 10643 4063
rect 10793 4029 10827 4063
rect 10885 4029 10919 4063
rect 12081 4029 12115 4063
rect 9137 3961 9171 3995
rect 9965 3961 9999 3995
rect 1869 3893 1903 3927
rect 8585 3893 8619 3927
rect 10793 3893 10827 3927
rect 7021 3689 7055 3723
rect 9873 3689 9907 3723
rect 10701 3689 10735 3723
rect 1593 3621 1627 3655
rect 6745 3553 6779 3587
rect 7297 3553 7331 3587
rect 9597 3553 9631 3587
rect 10149 3553 10183 3587
rect 11989 3553 12023 3587
rect 1409 3485 1443 3519
rect 7113 3485 7147 3519
rect 9965 3485 9999 3519
rect 10609 3485 10643 3519
rect 12265 3485 12299 3519
rect 6837 3417 6871 3451
rect 9689 3417 9723 3451
rect 8585 3145 8619 3179
rect 9689 3145 9723 3179
rect 12173 3145 12207 3179
rect 8493 3077 8527 3111
rect 12081 3077 12115 3111
rect 1409 3009 1443 3043
rect 8769 3009 8803 3043
rect 8953 3009 8987 3043
rect 10425 3009 10459 3043
rect 10701 3009 10735 3043
rect 8401 2941 8435 2975
rect 1593 2873 1627 2907
rect 4169 2601 4203 2635
rect 10793 2601 10827 2635
rect 11713 2601 11747 2635
rect 3801 2533 3835 2567
rect 6745 2533 6779 2567
rect 9321 2533 9355 2567
rect 1961 2397 1995 2431
rect 2881 2397 2915 2431
rect 3801 2397 3835 2431
rect 3985 2397 4019 2431
rect 5457 2397 5491 2431
rect 6561 2397 6595 2431
rect 7389 2397 7423 2431
rect 8033 2397 8067 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 10977 2397 11011 2431
rect 11621 2397 11655 2431
rect 1777 2329 1811 2363
rect 2697 2329 2731 2363
rect 5273 2329 5307 2363
rect 7849 2329 7883 2363
rect 7205 2261 7239 2295
rect 10149 2261 10183 2295
<< metal1 >>
rect 8018 13676 8024 13728
rect 8076 13716 8082 13728
rect 9766 13716 9772 13728
rect 8076 13688 9772 13716
rect 8076 13676 8082 13688
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 1104 13626 12972 13648
rect 1104 13574 2960 13626
rect 3012 13574 3024 13626
rect 3076 13574 3088 13626
rect 3140 13574 3152 13626
rect 3204 13574 6916 13626
rect 6968 13574 6980 13626
rect 7032 13574 7044 13626
rect 7096 13574 7108 13626
rect 7160 13574 10872 13626
rect 10924 13574 10936 13626
rect 10988 13574 11000 13626
rect 11052 13574 11064 13626
rect 11116 13574 12972 13626
rect 1104 13552 12972 13574
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 5408 13484 9352 13512
rect 5408 13472 5414 13484
rect 3418 13404 3424 13456
rect 3476 13444 3482 13456
rect 3476 13416 5212 13444
rect 3476 13404 3482 13416
rect 1762 13376 1768 13388
rect 1723 13348 1768 13376
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 1854 13336 1860 13388
rect 1912 13376 1918 13388
rect 1912 13348 3832 13376
rect 1912 13336 1918 13348
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 2774 13308 2780 13320
rect 2547 13280 2780 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 3804 13317 3832 13348
rect 3789 13311 3847 13317
rect 3789 13277 3801 13311
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 4430 13268 4436 13320
rect 4488 13308 4494 13320
rect 5184 13317 5212 13416
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 6733 13447 6791 13453
rect 6733 13444 6745 13447
rect 5776 13416 6745 13444
rect 5776 13404 5782 13416
rect 6733 13413 6745 13416
rect 6779 13413 6791 13447
rect 6733 13407 6791 13413
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 7469 13447 7527 13453
rect 7469 13444 7481 13447
rect 7340 13416 7481 13444
rect 7340 13404 7346 13416
rect 7469 13413 7481 13416
rect 7515 13413 7527 13447
rect 7469 13407 7527 13413
rect 9324 13444 9352 13484
rect 9324 13416 12204 13444
rect 4525 13311 4583 13317
rect 4525 13308 4537 13311
rect 4488 13280 4537 13308
rect 4488 13268 4494 13280
rect 4525 13277 4537 13280
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 5169 13311 5227 13317
rect 5169 13277 5181 13311
rect 5215 13277 5227 13311
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 5169 13271 5227 13277
rect 6886 13280 7665 13308
rect 1486 13200 1492 13252
rect 1544 13240 1550 13252
rect 1949 13243 2007 13249
rect 1949 13240 1961 13243
rect 1544 13212 1961 13240
rect 1544 13200 1550 13212
rect 1949 13209 1961 13212
rect 1995 13209 2007 13243
rect 1949 13203 2007 13209
rect 5442 13200 5448 13252
rect 5500 13240 5506 13252
rect 6886 13240 6914 13280
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 8294 13268 8300 13320
rect 8352 13308 8358 13320
rect 9324 13317 9352 13416
rect 10962 13376 10968 13388
rect 9508 13348 10824 13376
rect 10923 13348 10968 13376
rect 9508 13317 9536 13348
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8352 13280 8401 13308
rect 8352 13268 8358 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13277 9551 13311
rect 9493 13271 9551 13277
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 9824 13280 10701 13308
rect 9824 13268 9830 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10796 13308 10824 13348
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 12176 13385 12204 13416
rect 12161 13379 12219 13385
rect 11348 13348 12112 13376
rect 11348 13308 11376 13348
rect 10796 13280 11376 13308
rect 11701 13311 11759 13317
rect 10689 13271 10747 13277
rect 11701 13277 11713 13311
rect 11747 13277 11759 13311
rect 11882 13308 11888 13320
rect 11843 13280 11888 13308
rect 11701 13271 11759 13277
rect 5500 13212 6914 13240
rect 6953 13243 7011 13249
rect 5500 13200 5506 13212
rect 6953 13209 6965 13243
rect 6999 13240 7011 13243
rect 9582 13240 9588 13252
rect 6999 13212 9588 13240
rect 6999 13209 7011 13212
rect 6953 13203 7011 13209
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 11716 13240 11744 13271
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 12084 13252 12112 13348
rect 12161 13345 12173 13379
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 9723 13212 11744 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 12066 13249 12072 13252
rect 12023 13243 12072 13249
rect 11848 13212 11893 13240
rect 11848 13200 11854 13212
rect 12023 13209 12035 13243
rect 12069 13209 12072 13243
rect 12023 13203 12072 13209
rect 12066 13200 12072 13203
rect 12124 13200 12130 13252
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3973 13175 4031 13181
rect 3973 13141 3985 13175
rect 4019 13172 4031 13175
rect 4522 13172 4528 13184
rect 4019 13144 4528 13172
rect 4019 13141 4031 13144
rect 3973 13135 4031 13141
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 4709 13175 4767 13181
rect 4709 13141 4721 13175
rect 4755 13172 4767 13175
rect 5258 13172 5264 13184
rect 4755 13144 5264 13172
rect 4755 13141 4767 13144
rect 4709 13135 4767 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5353 13175 5411 13181
rect 5353 13141 5365 13175
rect 5399 13172 5411 13175
rect 6546 13172 6552 13184
rect 5399 13144 6552 13172
rect 5399 13141 5411 13144
rect 5353 13135 5411 13141
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 7524 13144 8217 13172
rect 7524 13132 7530 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 8205 13135 8263 13141
rect 8294 13132 8300 13184
rect 8352 13172 8358 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 8352 13144 11529 13172
rect 8352 13132 8358 13144
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 1104 13082 12972 13104
rect 1104 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 8894 13082
rect 8946 13030 8958 13082
rect 9010 13030 9022 13082
rect 9074 13030 9086 13082
rect 9138 13030 12972 13082
rect 1104 13008 12972 13030
rect 2682 12928 2688 12980
rect 2740 12968 2746 12980
rect 9858 12968 9864 12980
rect 2740 12940 9864 12968
rect 2740 12928 2746 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 11701 12971 11759 12977
rect 11701 12937 11713 12971
rect 11747 12968 11759 12971
rect 11790 12968 11796 12980
rect 11747 12940 11796 12968
rect 11747 12937 11759 12940
rect 11701 12931 11759 12937
rect 11790 12928 11796 12940
rect 11848 12968 11854 12980
rect 11974 12968 11980 12980
rect 11848 12940 11980 12968
rect 11848 12928 11854 12940
rect 11974 12928 11980 12940
rect 12032 12928 12038 12980
rect 566 12860 572 12912
rect 624 12900 630 12912
rect 1765 12903 1823 12909
rect 1765 12900 1777 12903
rect 624 12872 1777 12900
rect 624 12860 630 12872
rect 1765 12869 1777 12872
rect 1811 12869 1823 12903
rect 1765 12863 1823 12869
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12900 2007 12903
rect 1995 12872 3924 12900
rect 1995 12869 2007 12872
rect 1949 12863 2007 12869
rect 3418 12832 3424 12844
rect 3379 12804 3424 12832
rect 3418 12792 3424 12804
rect 3476 12792 3482 12844
rect 3896 12832 3924 12872
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 4614 12900 4620 12912
rect 4028 12872 4073 12900
rect 4172 12872 4620 12900
rect 4028 12860 4034 12872
rect 4172 12832 4200 12872
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 5534 12860 5540 12912
rect 5592 12900 5598 12912
rect 9950 12900 9956 12912
rect 5592 12872 7328 12900
rect 5592 12860 5598 12872
rect 3896 12804 4200 12832
rect 4248 12835 4306 12841
rect 4248 12801 4260 12835
rect 4294 12832 4306 12835
rect 4338 12832 4344 12844
rect 4294 12804 4344 12832
rect 4294 12801 4306 12804
rect 4248 12795 4306 12801
rect 4338 12792 4344 12804
rect 4396 12792 4402 12844
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 7193 12835 7251 12841
rect 7193 12832 7205 12835
rect 4764 12804 7205 12832
rect 4764 12792 4770 12804
rect 7193 12801 7205 12804
rect 7239 12801 7251 12835
rect 7193 12795 7251 12801
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4430 12764 4436 12776
rect 3927 12736 4436 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 7101 12767 7159 12773
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7300 12764 7328 12872
rect 9048 12872 9956 12900
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 8294 12832 8300 12844
rect 7699 12804 8300 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 9048 12841 9076 12872
rect 9950 12860 9956 12872
rect 10008 12860 10014 12912
rect 10873 12903 10931 12909
rect 10873 12869 10885 12903
rect 10919 12900 10931 12903
rect 12158 12900 12164 12912
rect 10919 12872 12164 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9306 12832 9312 12844
rect 9267 12804 9312 12832
rect 9033 12795 9091 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 9766 12832 9772 12844
rect 9447 12804 9772 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 11698 12792 11704 12804
rect 11756 12832 11762 12844
rect 11882 12832 11888 12844
rect 11756 12804 11888 12832
rect 11756 12792 11762 12804
rect 11882 12792 11888 12804
rect 11940 12832 11946 12844
rect 11940 12804 12204 12832
rect 11940 12792 11946 12804
rect 12176 12773 12204 12804
rect 12161 12767 12219 12773
rect 7147 12736 11560 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 3329 12699 3387 12705
rect 3329 12665 3341 12699
rect 3375 12696 3387 12699
rect 4246 12696 4252 12708
rect 3375 12668 4252 12696
rect 3375 12665 3387 12668
rect 3329 12659 3387 12665
rect 4246 12656 4252 12668
rect 4304 12656 4310 12708
rect 6932 12696 6960 12727
rect 7282 12696 7288 12708
rect 6932 12668 7288 12696
rect 7282 12656 7288 12668
rect 7340 12656 7346 12708
rect 7558 12696 7564 12708
rect 7519 12668 7564 12696
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 9125 12699 9183 12705
rect 9125 12665 9137 12699
rect 9171 12696 9183 12699
rect 10318 12696 10324 12708
rect 9171 12668 10324 12696
rect 9171 12665 9183 12668
rect 9125 12659 9183 12665
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 10410 12656 10416 12708
rect 10468 12696 10474 12708
rect 11532 12705 11560 12736
rect 12161 12733 12173 12767
rect 12207 12733 12219 12767
rect 12161 12727 12219 12733
rect 10597 12699 10655 12705
rect 10597 12696 10609 12699
rect 10468 12668 10609 12696
rect 10468 12656 10474 12668
rect 10597 12665 10609 12668
rect 10643 12665 10655 12699
rect 10597 12659 10655 12665
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12665 11575 12699
rect 11517 12659 11575 12665
rect 4154 12628 4160 12640
rect 4115 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 10502 12628 10508 12640
rect 9631 12600 10508 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12069 12631 12127 12637
rect 12069 12628 12081 12631
rect 12032 12600 12081 12628
rect 12032 12588 12038 12600
rect 12069 12597 12081 12600
rect 12115 12597 12127 12631
rect 12069 12591 12127 12597
rect 1104 12538 12972 12560
rect 1104 12486 2960 12538
rect 3012 12486 3024 12538
rect 3076 12486 3088 12538
rect 3140 12486 3152 12538
rect 3204 12486 6916 12538
rect 6968 12486 6980 12538
rect 7032 12486 7044 12538
rect 7096 12486 7108 12538
rect 7160 12486 10872 12538
rect 10924 12486 10936 12538
rect 10988 12486 11000 12538
rect 11052 12486 11064 12538
rect 11116 12486 12972 12538
rect 1104 12464 12972 12486
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 3936 12396 4200 12424
rect 3936 12384 3942 12396
rect 3694 12316 3700 12368
rect 3752 12356 3758 12368
rect 4065 12359 4123 12365
rect 4065 12356 4077 12359
rect 3752 12328 4077 12356
rect 3752 12316 3758 12328
rect 4065 12325 4077 12328
rect 4111 12325 4123 12359
rect 4172 12356 4200 12396
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 10873 12427 10931 12433
rect 10873 12424 10885 12427
rect 10652 12396 10885 12424
rect 10652 12384 10658 12396
rect 10873 12393 10885 12396
rect 10919 12393 10931 12427
rect 10873 12387 10931 12393
rect 10778 12356 10784 12368
rect 4172 12328 10784 12356
rect 4065 12319 4123 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 4154 12288 4160 12300
rect 2746 12260 4160 12288
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 2746 12220 2774 12260
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 8386 12288 8392 12300
rect 4263 12260 8392 12288
rect 3786 12220 3792 12232
rect 1719 12192 2774 12220
rect 3747 12192 3792 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 1412 12152 1440 12183
rect 3786 12180 3792 12192
rect 3844 12180 3850 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3896 12192 3985 12220
rect 1762 12152 1768 12164
rect 1412 12124 1768 12152
rect 1762 12112 1768 12124
rect 1820 12112 1826 12164
rect 2406 12084 2412 12096
rect 2367 12056 2412 12084
rect 2406 12044 2412 12056
rect 2464 12044 2470 12096
rect 3896 12084 3924 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 4263 12220 4291 12260
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 9490 12248 9496 12300
rect 9548 12288 9554 12300
rect 11977 12291 12035 12297
rect 11977 12288 11989 12291
rect 9548 12260 11989 12288
rect 9548 12248 9554 12260
rect 11977 12257 11989 12260
rect 12023 12257 12035 12291
rect 11977 12251 12035 12257
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 13446 12288 13452 12300
rect 12299 12260 13452 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 13446 12248 13452 12260
rect 13504 12248 13510 12300
rect 4120 12192 4291 12220
rect 4120 12180 4126 12192
rect 4338 12180 4344 12232
rect 4396 12220 4402 12232
rect 5994 12220 6000 12232
rect 4396 12192 6000 12220
rect 4396 12180 4402 12192
rect 5994 12180 6000 12192
rect 6052 12180 6058 12232
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9272 12192 9873 12220
rect 9272 12180 9278 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 4430 12112 4436 12164
rect 4488 12152 4494 12164
rect 4488 12124 9996 12152
rect 4488 12112 4494 12124
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 3896 12056 4261 12084
rect 4249 12053 4261 12056
rect 4295 12084 4307 12087
rect 5810 12084 5816 12096
rect 4295 12056 5816 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 7708 12056 9689 12084
rect 7708 12044 7714 12056
rect 9677 12053 9689 12056
rect 9723 12053 9735 12087
rect 9968 12084 9996 12124
rect 10042 12112 10048 12164
rect 10100 12152 10106 12164
rect 10781 12155 10839 12161
rect 10781 12152 10793 12155
rect 10100 12124 10793 12152
rect 10100 12112 10106 12124
rect 10781 12121 10793 12124
rect 10827 12121 10839 12155
rect 10781 12115 10839 12121
rect 12066 12084 12072 12096
rect 9968 12056 12072 12084
rect 9677 12047 9735 12053
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 1104 11994 12972 12016
rect 1104 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 8894 11994
rect 8946 11942 8958 11994
rect 9010 11942 9022 11994
rect 9074 11942 9086 11994
rect 9138 11942 12972 11994
rect 1104 11920 12972 11942
rect 3237 11883 3295 11889
rect 3237 11849 3249 11883
rect 3283 11880 3295 11883
rect 9306 11880 9312 11892
rect 3283 11852 9312 11880
rect 3283 11849 3295 11852
rect 3237 11843 3295 11849
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3252 11744 3280 11843
rect 9306 11840 9312 11852
rect 9364 11880 9370 11892
rect 12253 11883 12311 11889
rect 12253 11880 12265 11883
rect 9364 11852 12265 11880
rect 9364 11840 9370 11852
rect 12253 11849 12265 11852
rect 12299 11849 12311 11883
rect 12253 11843 12311 11849
rect 9674 11812 9680 11824
rect 3344 11784 9680 11812
rect 3344 11753 3372 11784
rect 9674 11772 9680 11784
rect 9732 11772 9738 11824
rect 9784 11784 12020 11812
rect 3007 11716 3280 11744
rect 3329 11747 3387 11753
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3329 11713 3341 11747
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 1394 11676 1400 11688
rect 1355 11648 1400 11676
rect 1394 11636 1400 11648
rect 1452 11636 1458 11688
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11645 1731 11679
rect 1673 11639 1731 11645
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 3344 11676 3372 11707
rect 6362 11704 6368 11756
rect 6420 11744 6426 11756
rect 6532 11747 6590 11753
rect 6532 11744 6544 11747
rect 6420 11716 6544 11744
rect 6420 11704 6426 11716
rect 6532 11713 6544 11716
rect 6578 11713 6590 11747
rect 6671 11747 6729 11753
rect 6671 11744 6683 11747
rect 6532 11707 6590 11713
rect 6657 11713 6683 11744
rect 6717 11713 6729 11747
rect 6914 11744 6920 11756
rect 6827 11716 6920 11744
rect 6657 11707 6729 11713
rect 2823 11648 3372 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 1688 11540 1716 11639
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 6657 11676 6685 11707
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 8294 11744 8300 11756
rect 6972 11716 8300 11744
rect 6972 11704 6978 11716
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 8386 11704 8392 11756
rect 8444 11744 8450 11756
rect 9784 11744 9812 11784
rect 8444 11716 9812 11744
rect 10321 11747 10379 11753
rect 8444 11704 8450 11716
rect 10321 11713 10333 11747
rect 10367 11744 10379 11747
rect 10686 11744 10692 11756
rect 10367 11716 10692 11744
rect 10367 11713 10379 11716
rect 10321 11707 10379 11713
rect 10686 11704 10692 11716
rect 10744 11704 10750 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 11698 11744 11704 11756
rect 10836 11716 10881 11744
rect 11659 11716 11704 11744
rect 10836 11704 10842 11716
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11992 11753 12020 11784
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12066 11704 12072 11756
rect 12124 11744 12130 11756
rect 12124 11716 12169 11744
rect 12124 11704 12130 11716
rect 5776 11648 6685 11676
rect 5776 11636 5782 11648
rect 8018 11636 8024 11688
rect 8076 11676 8082 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 8076 11648 11805 11676
rect 8076 11636 8082 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 3053 11611 3111 11617
rect 3053 11577 3065 11611
rect 3099 11608 3111 11611
rect 6454 11608 6460 11620
rect 3099 11580 6460 11608
rect 3099 11577 3111 11580
rect 3053 11571 3111 11577
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 10873 11611 10931 11617
rect 10873 11608 10885 11611
rect 9508 11580 10885 11608
rect 3602 11540 3608 11552
rect 1688 11512 3608 11540
rect 3602 11500 3608 11512
rect 3660 11540 3666 11552
rect 3878 11540 3884 11552
rect 3660 11512 3884 11540
rect 3660 11500 3666 11512
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 4028 11512 6377 11540
rect 4028 11500 4034 11512
rect 6365 11509 6377 11512
rect 6411 11509 6423 11543
rect 6365 11503 6423 11509
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 9214 11500 9220 11552
rect 9272 11540 9278 11552
rect 9508 11540 9536 11580
rect 10873 11577 10885 11580
rect 10919 11577 10931 11611
rect 10873 11571 10931 11577
rect 9272 11512 9536 11540
rect 9272 11500 9278 11512
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 10137 11543 10195 11549
rect 10137 11540 10149 11543
rect 9824 11512 10149 11540
rect 9824 11500 9830 11512
rect 10137 11509 10149 11512
rect 10183 11509 10195 11543
rect 10137 11503 10195 11509
rect 1104 11450 12972 11472
rect 1104 11398 2960 11450
rect 3012 11398 3024 11450
rect 3076 11398 3088 11450
rect 3140 11398 3152 11450
rect 3204 11398 6916 11450
rect 6968 11398 6980 11450
rect 7032 11398 7044 11450
rect 7096 11398 7108 11450
rect 7160 11398 10872 11450
rect 10924 11398 10936 11450
rect 10988 11398 11000 11450
rect 11052 11398 11064 11450
rect 11116 11398 12972 11450
rect 1104 11376 12972 11398
rect 4706 11336 4712 11348
rect 4667 11308 4712 11336
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 5721 11339 5779 11345
rect 5721 11305 5733 11339
rect 5767 11336 5779 11339
rect 9766 11336 9772 11348
rect 5767 11308 9772 11336
rect 5767 11305 5779 11308
rect 5721 11299 5779 11305
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 12069 11339 12127 11345
rect 12069 11336 12081 11339
rect 10284 11308 12081 11336
rect 10284 11296 10290 11308
rect 12069 11305 12081 11308
rect 12115 11305 12127 11339
rect 12069 11299 12127 11305
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 9214 11268 9220 11280
rect 3936 11240 9220 11268
rect 3936 11228 3942 11240
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 5258 11200 5264 11212
rect 4764 11172 5264 11200
rect 4764 11160 4770 11172
rect 5258 11160 5264 11172
rect 5316 11160 5322 11212
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 4062 11132 4068 11144
rect 3476 11104 4068 11132
rect 3476 11092 3482 11104
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 5828 11141 5856 11240
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 11333 11271 11391 11277
rect 11333 11268 11345 11271
rect 9364 11240 11345 11268
rect 9364 11228 9370 11240
rect 11333 11237 11345 11240
rect 11379 11237 11391 11271
rect 11333 11231 11391 11237
rect 5905 11203 5963 11209
rect 5905 11169 5917 11203
rect 5951 11169 5963 11203
rect 7558 11200 7564 11212
rect 5905 11163 5963 11169
rect 6104 11172 7564 11200
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11132 4859 11135
rect 5721 11135 5779 11141
rect 5721 11132 5733 11135
rect 4847 11104 5733 11132
rect 4847 11101 4859 11104
rect 4801 11095 4859 11101
rect 5721 11101 5733 11104
rect 5767 11101 5779 11135
rect 5721 11095 5779 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 3786 11024 3792 11076
rect 3844 11064 3850 11076
rect 5920 11064 5948 11163
rect 6104 11141 6132 11172
rect 7558 11160 7564 11172
rect 7616 11200 7622 11212
rect 11146 11200 11152 11212
rect 7616 11172 11152 11200
rect 7616 11160 7622 11172
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11609 11203 11667 11209
rect 11609 11200 11621 11203
rect 11256 11172 11621 11200
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11101 6147 11135
rect 6089 11095 6147 11101
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6196 11064 6224 11095
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 10594 11132 10600 11144
rect 6512 11104 10600 11132
rect 6512 11092 6518 11104
rect 10594 11092 10600 11104
rect 10652 11092 10658 11144
rect 11057 11135 11115 11141
rect 11057 11101 11069 11135
rect 11103 11132 11115 11135
rect 11256 11132 11284 11172
rect 11609 11169 11621 11172
rect 11655 11169 11667 11203
rect 11609 11163 11667 11169
rect 11103 11104 11284 11132
rect 11425 11135 11483 11141
rect 11103 11101 11115 11104
rect 11057 11095 11115 11101
rect 11425 11101 11437 11135
rect 11471 11101 11483 11135
rect 12250 11132 12256 11144
rect 12211 11104 12256 11132
rect 11425 11095 11483 11101
rect 6365 11067 6423 11073
rect 3844 11036 5948 11064
rect 6012 11036 6316 11064
rect 3844 11024 3850 11036
rect 5258 10956 5264 11008
rect 5316 10996 5322 11008
rect 6012 10996 6040 11036
rect 5316 10968 6040 10996
rect 6288 10996 6316 11036
rect 6365 11033 6377 11067
rect 6411 11064 6423 11067
rect 7282 11064 7288 11076
rect 6411 11036 7288 11064
rect 6411 11033 6423 11036
rect 6365 11027 6423 11033
rect 7282 11024 7288 11036
rect 7340 11024 7346 11076
rect 7392 11036 8156 11064
rect 7392 10996 7420 11036
rect 6288 10968 7420 10996
rect 8128 10996 8156 11036
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 10226 11064 10232 11076
rect 8260 11036 10232 11064
rect 8260 11024 8266 11036
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 11072 11064 11100 11095
rect 10336 11036 11100 11064
rect 10336 10996 10364 11036
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11440 11064 11468 11095
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 11204 11036 11468 11064
rect 11204 11024 11210 11036
rect 8128 10968 10364 10996
rect 5316 10956 5322 10968
rect 10410 10956 10416 11008
rect 10468 10996 10474 11008
rect 10686 10996 10692 11008
rect 10468 10968 10692 10996
rect 10468 10956 10474 10968
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 1104 10906 12972 10928
rect 1104 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 8894 10906
rect 8946 10854 8958 10906
rect 9010 10854 9022 10906
rect 9074 10854 9086 10906
rect 9138 10854 12972 10906
rect 1104 10832 12972 10854
rect 4249 10795 4307 10801
rect 4249 10761 4261 10795
rect 4295 10792 4307 10795
rect 5534 10792 5540 10804
rect 4295 10764 5540 10792
rect 4295 10761 4307 10764
rect 4249 10755 4307 10761
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10656 4031 10659
rect 4264 10656 4292 10755
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 9398 10792 9404 10804
rect 6420 10764 9404 10792
rect 6420 10752 6426 10764
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 4706 10684 4712 10736
rect 4764 10724 4770 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4764 10696 5089 10724
rect 4764 10684 4770 10696
rect 5077 10693 5089 10696
rect 5123 10693 5135 10727
rect 5077 10687 5135 10693
rect 5169 10727 5227 10733
rect 5169 10693 5181 10727
rect 5215 10724 5227 10727
rect 7742 10724 7748 10736
rect 5215 10696 7748 10724
rect 5215 10693 5227 10696
rect 5169 10687 5227 10693
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 4019 10628 4292 10656
rect 4985 10659 5043 10665
rect 4019 10625 4031 10628
rect 3973 10619 4031 10625
rect 4985 10625 4997 10659
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 11790 10656 11796 10668
rect 5399 10628 11796 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10588 3847 10591
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 3835 10560 4353 10588
rect 3835 10557 3847 10560
rect 3789 10551 3847 10557
rect 3988 10452 4016 10560
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 5000 10588 5028 10619
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 8662 10588 8668 10600
rect 5000 10560 8668 10588
rect 4341 10551 4399 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 4065 10523 4123 10529
rect 4065 10489 4077 10523
rect 4111 10520 4123 10523
rect 6178 10520 6184 10532
rect 4111 10492 6184 10520
rect 4111 10489 4123 10492
rect 4065 10483 4123 10489
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 11882 10520 11888 10532
rect 6328 10492 11888 10520
rect 6328 10480 6334 10492
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 4801 10455 4859 10461
rect 4801 10452 4813 10455
rect 3988 10424 4813 10452
rect 4801 10421 4813 10424
rect 4847 10452 4859 10455
rect 7374 10452 7380 10464
rect 4847 10424 7380 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 7374 10412 7380 10424
rect 7432 10452 7438 10464
rect 7558 10452 7564 10464
rect 7432 10424 7564 10452
rect 7432 10412 7438 10424
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 1104 10362 12972 10384
rect 1104 10310 2960 10362
rect 3012 10310 3024 10362
rect 3076 10310 3088 10362
rect 3140 10310 3152 10362
rect 3204 10310 6916 10362
rect 6968 10310 6980 10362
rect 7032 10310 7044 10362
rect 7096 10310 7108 10362
rect 7160 10310 10872 10362
rect 10924 10310 10936 10362
rect 10988 10310 11000 10362
rect 11052 10310 11064 10362
rect 11116 10310 12972 10362
rect 1104 10288 12972 10310
rect 2593 10251 2651 10257
rect 2593 10217 2605 10251
rect 2639 10248 2651 10251
rect 3786 10248 3792 10260
rect 2639 10220 3792 10248
rect 2639 10217 2651 10220
rect 2593 10211 2651 10217
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 7466 10248 7472 10260
rect 4396 10220 7472 10248
rect 4396 10208 4402 10220
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 10008 10220 10057 10248
rect 10008 10208 10014 10220
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10045 10211 10103 10217
rect 12069 10251 12127 10257
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 12158 10248 12164 10260
rect 12115 10220 12164 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 3326 10140 3332 10192
rect 3384 10180 3390 10192
rect 8665 10183 8723 10189
rect 8665 10180 8677 10183
rect 3384 10152 8677 10180
rect 3384 10140 3390 10152
rect 8665 10149 8677 10152
rect 8711 10149 8723 10183
rect 8665 10143 8723 10149
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 9490 10180 9496 10192
rect 8803 10152 9496 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 5920 10084 9260 10112
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 4338 10044 4344 10056
rect 2731 10016 4344 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4522 10004 4528 10056
rect 4580 10044 4586 10056
rect 5920 10044 5948 10084
rect 9232 10053 9260 10084
rect 9324 10053 9352 10152
rect 9490 10140 9496 10152
rect 9548 10140 9554 10192
rect 4580 10016 5948 10044
rect 8665 10047 8723 10053
rect 4580 10004 4586 10016
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8711 10016 8953 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9309 10047 9367 10053
rect 9309 10013 9321 10047
rect 9355 10013 9367 10047
rect 9309 10007 9367 10013
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 9953 10047 10011 10053
rect 9953 10044 9965 10047
rect 9916 10016 9965 10044
rect 9916 10004 9922 10016
rect 9953 10013 9965 10016
rect 9999 10013 10011 10047
rect 10962 10044 10968 10056
rect 10923 10016 10968 10044
rect 9953 10007 10011 10013
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 12250 10044 12256 10056
rect 12211 10016 12256 10044
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 1854 9976 1860 9988
rect 1815 9948 1860 9976
rect 1854 9936 1860 9948
rect 1912 9936 1918 9988
rect 9125 9979 9183 9985
rect 9125 9976 9137 9979
rect 4448 9948 9137 9976
rect 1946 9908 1952 9920
rect 1907 9880 1952 9908
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4448 9917 4476 9948
rect 9125 9945 9137 9948
rect 9171 9945 9183 9979
rect 9125 9939 9183 9945
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4120 9880 4445 9908
rect 4120 9868 4126 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4433 9871 4491 9877
rect 5534 9868 5540 9920
rect 5592 9908 5598 9920
rect 8665 9911 8723 9917
rect 8665 9908 8677 9911
rect 5592 9880 8677 9908
rect 5592 9868 5598 9880
rect 8665 9877 8677 9880
rect 8711 9877 8723 9911
rect 8665 9871 8723 9877
rect 8754 9868 8760 9920
rect 8812 9908 8818 9920
rect 9493 9911 9551 9917
rect 9493 9908 9505 9911
rect 8812 9880 9505 9908
rect 8812 9868 8818 9880
rect 9493 9877 9505 9880
rect 9539 9877 9551 9911
rect 9493 9871 9551 9877
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 11057 9911 11115 9917
rect 11057 9908 11069 9911
rect 10284 9880 11069 9908
rect 10284 9868 10290 9880
rect 11057 9877 11069 9880
rect 11103 9877 11115 9911
rect 11057 9871 11115 9877
rect 1104 9818 12972 9840
rect 1104 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 8894 9818
rect 8946 9766 8958 9818
rect 9010 9766 9022 9818
rect 9074 9766 9086 9818
rect 9138 9766 12972 9818
rect 1104 9744 12972 9766
rect 1946 9664 1952 9716
rect 2004 9704 2010 9716
rect 6270 9704 6276 9716
rect 2004 9676 6276 9704
rect 2004 9664 2010 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 6362 9664 6368 9716
rect 6420 9704 6426 9716
rect 10962 9704 10968 9716
rect 6420 9676 10968 9704
rect 6420 9664 6426 9676
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11514 9636 11520 9648
rect 8312 9608 11520 9636
rect 6638 9568 6644 9580
rect 6599 9540 6644 9568
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 8312 9577 8340 9608
rect 11514 9596 11520 9608
rect 11572 9596 11578 9648
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9537 8355 9571
rect 9306 9568 9312 9580
rect 9267 9540 9312 9568
rect 8297 9531 8355 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9033 9503 9091 9509
rect 9033 9500 9045 9503
rect 8619 9472 9045 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 9033 9469 9045 9472
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9048 9432 9076 9463
rect 10042 9432 10048 9444
rect 9048 9404 9168 9432
rect 10003 9404 10048 9432
rect 6730 9364 6736 9376
rect 6691 9336 6736 9364
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7432 9336 7573 9364
rect 7432 9324 7438 9336
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 9140 9364 9168 9404
rect 10042 9392 10048 9404
rect 10100 9392 10106 9444
rect 9306 9364 9312 9376
rect 9140 9336 9312 9364
rect 7561 9327 7619 9333
rect 9306 9324 9312 9336
rect 9364 9364 9370 9376
rect 10686 9364 10692 9376
rect 9364 9336 10692 9364
rect 9364 9324 9370 9336
rect 10686 9324 10692 9336
rect 10744 9364 10750 9376
rect 11238 9364 11244 9376
rect 10744 9336 11244 9364
rect 10744 9324 10750 9336
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 1104 9274 12972 9296
rect 1104 9222 2960 9274
rect 3012 9222 3024 9274
rect 3076 9222 3088 9274
rect 3140 9222 3152 9274
rect 3204 9222 6916 9274
rect 6968 9222 6980 9274
rect 7032 9222 7044 9274
rect 7096 9222 7108 9274
rect 7160 9222 10872 9274
rect 10924 9222 10936 9274
rect 10988 9222 11000 9274
rect 11052 9222 11064 9274
rect 11116 9222 12972 9274
rect 1104 9200 12972 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 5077 9163 5135 9169
rect 2915 9132 5028 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 5000 9092 5028 9132
rect 5077 9129 5089 9163
rect 5123 9160 5135 9163
rect 5442 9160 5448 9172
rect 5123 9132 5448 9160
rect 5123 9129 5135 9132
rect 5077 9123 5135 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 9582 9160 9588 9172
rect 6696 9132 9588 9160
rect 6696 9120 6702 9132
rect 9582 9120 9588 9132
rect 9640 9120 9646 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 9769 9163 9827 9169
rect 9769 9160 9781 9163
rect 9732 9132 9781 9160
rect 9732 9120 9738 9132
rect 9769 9129 9781 9132
rect 9815 9129 9827 9163
rect 11330 9160 11336 9172
rect 9769 9123 9827 9129
rect 9876 9132 11336 9160
rect 9876 9092 9904 9132
rect 11330 9120 11336 9132
rect 11388 9120 11394 9172
rect 5000 9064 9904 9092
rect 9950 9052 9956 9104
rect 10008 9052 10014 9104
rect 1762 8984 1768 9036
rect 1820 9024 1826 9036
rect 1857 9027 1915 9033
rect 1857 9024 1869 9027
rect 1820 8996 1869 9024
rect 1820 8984 1826 8996
rect 1857 8993 1869 8996
rect 1903 8993 1915 9027
rect 1857 8987 1915 8993
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 9024 6055 9027
rect 8478 9024 8484 9036
rect 6043 8996 8484 9024
rect 6043 8993 6055 8996
rect 5997 8987 6055 8993
rect 1872 8888 1900 8987
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 9968 9024 9996 9052
rect 9968 8996 10180 9024
rect 2130 8956 2136 8968
rect 2091 8928 2136 8956
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 2746 8928 4077 8956
rect 2746 8900 2774 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 5626 8956 5632 8968
rect 4387 8928 5632 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 5721 8959 5779 8965
rect 5721 8925 5733 8959
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 2746 8888 2780 8900
rect 1872 8860 2780 8888
rect 2774 8848 2780 8860
rect 2832 8848 2838 8900
rect 5736 8888 5764 8919
rect 5810 8916 5816 8968
rect 5868 8956 5874 8968
rect 6089 8959 6147 8965
rect 5868 8928 5913 8956
rect 5868 8916 5874 8928
rect 6089 8925 6101 8959
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 5994 8888 6000 8900
rect 5736 8860 6000 8888
rect 5994 8848 6000 8860
rect 6052 8848 6058 8900
rect 5534 8820 5540 8832
rect 5495 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 6104 8820 6132 8919
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 10152 8965 10180 8996
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 6604 8928 9965 8956
rect 6604 8916 6610 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 10137 8919 10195 8925
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 9674 8888 9680 8900
rect 6788 8860 9680 8888
rect 6788 8848 6794 8860
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10045 8891 10103 8897
rect 10045 8888 10057 8891
rect 9916 8860 10057 8888
rect 9916 8848 9922 8860
rect 10045 8857 10057 8860
rect 10091 8857 10103 8891
rect 10045 8851 10103 8857
rect 11606 8820 11612 8832
rect 6104 8792 11612 8820
rect 11606 8780 11612 8792
rect 11664 8780 11670 8832
rect 1104 8730 12972 8752
rect 1104 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8894 8730
rect 8946 8678 8958 8730
rect 9010 8678 9022 8730
rect 9074 8678 9086 8730
rect 9138 8678 12972 8730
rect 1104 8656 12972 8678
rect 2130 8576 2136 8628
rect 2188 8616 2194 8628
rect 2188 8588 2774 8616
rect 2188 8576 2194 8588
rect 2746 8412 2774 8588
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9732 8588 9996 8616
rect 9732 8576 9738 8588
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 9769 8551 9827 8557
rect 9769 8548 9781 8551
rect 8352 8520 9781 8548
rect 8352 8508 8358 8520
rect 9769 8517 9781 8520
rect 9815 8517 9827 8551
rect 9769 8511 9827 8517
rect 8665 8483 8723 8489
rect 8665 8449 8677 8483
rect 8711 8480 8723 8483
rect 9582 8480 9588 8492
rect 8711 8452 9444 8480
rect 9543 8452 9588 8480
rect 8711 8449 8723 8452
rect 8665 8443 8723 8449
rect 8941 8415 8999 8421
rect 2746 8384 8340 8412
rect 7929 8347 7987 8353
rect 7929 8313 7941 8347
rect 7975 8344 7987 8347
rect 8110 8344 8116 8356
rect 7975 8316 8116 8344
rect 7975 8313 7987 8316
rect 7929 8307 7987 8313
rect 8110 8304 8116 8316
rect 8168 8304 8174 8356
rect 8312 8276 8340 8384
rect 8941 8381 8953 8415
rect 8987 8412 8999 8415
rect 9306 8412 9312 8424
rect 8987 8384 9312 8412
rect 8987 8381 8999 8384
rect 8941 8375 8999 8381
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 9416 8412 9444 8452
rect 9582 8440 9588 8452
rect 9640 8440 9646 8492
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 9968 8489 9996 8588
rect 9953 8483 10011 8489
rect 9732 8452 9777 8480
rect 9732 8440 9738 8452
rect 9953 8449 9965 8483
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 10686 8412 10692 8424
rect 9416 8384 10692 8412
rect 10686 8372 10692 8384
rect 10744 8372 10750 8424
rect 9398 8344 9404 8356
rect 9359 8316 9404 8344
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 9858 8344 9864 8356
rect 9508 8316 9864 8344
rect 9508 8276 9536 8316
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 8312 8248 9536 8276
rect 1104 8186 12972 8208
rect 1104 8134 2960 8186
rect 3012 8134 3024 8186
rect 3076 8134 3088 8186
rect 3140 8134 3152 8186
rect 3204 8134 6916 8186
rect 6968 8134 6980 8186
rect 7032 8134 7044 8186
rect 7096 8134 7108 8186
rect 7160 8134 10872 8186
rect 10924 8134 10936 8186
rect 10988 8134 11000 8186
rect 11052 8134 11064 8186
rect 11116 8134 12972 8186
rect 1104 8112 12972 8134
rect 3326 8072 3332 8084
rect 2884 8044 3332 8072
rect 2884 8016 2912 8044
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 2590 8004 2596 8016
rect 1596 7976 2596 8004
rect 1596 7877 1624 7976
rect 2590 7964 2596 7976
rect 2648 7964 2654 8016
rect 2866 7964 2872 8016
rect 2924 7964 2930 8016
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7834 8004 7840 8016
rect 6788 7976 7840 8004
rect 6788 7964 6794 7976
rect 7834 7964 7840 7976
rect 7892 7964 7898 8016
rect 2133 7939 2191 7945
rect 2133 7905 2145 7939
rect 2179 7936 2191 7939
rect 2685 7939 2743 7945
rect 2685 7936 2697 7939
rect 2179 7908 2697 7936
rect 2179 7905 2191 7908
rect 2133 7899 2191 7905
rect 2685 7905 2697 7908
rect 2731 7936 2743 7939
rect 3234 7936 3240 7948
rect 2731 7908 3240 7936
rect 2731 7905 2743 7908
rect 2685 7899 2743 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 11974 7936 11980 7948
rect 11935 7908 11980 7936
rect 11974 7896 11980 7908
rect 12032 7896 12038 7948
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7837 1639 7871
rect 1581 7831 1639 7837
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2332 7800 2360 7831
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 7834 7868 7840 7880
rect 3568 7840 7840 7868
rect 3568 7828 3574 7840
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 12250 7868 12256 7880
rect 12211 7840 12256 7868
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 2593 7803 2651 7809
rect 2593 7800 2605 7803
rect 2332 7772 2605 7800
rect 2593 7769 2605 7772
rect 2639 7769 2651 7803
rect 2593 7763 2651 7769
rect 1486 7732 1492 7744
rect 1447 7704 1492 7732
rect 1486 7692 1492 7704
rect 1544 7692 1550 7744
rect 2498 7732 2504 7744
rect 2459 7704 2504 7732
rect 2498 7692 2504 7704
rect 2556 7692 2562 7744
rect 2608 7732 2636 7763
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 9674 7800 9680 7812
rect 2740 7772 9680 7800
rect 2740 7760 2746 7772
rect 9674 7760 9680 7772
rect 9732 7760 9738 7812
rect 3510 7732 3516 7744
rect 2608 7704 3516 7732
rect 3510 7692 3516 7704
rect 3568 7732 3574 7744
rect 3970 7732 3976 7744
rect 3568 7704 3976 7732
rect 3568 7692 3574 7704
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 8018 7732 8024 7744
rect 6512 7704 8024 7732
rect 6512 7692 6518 7704
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 1104 7642 12972 7664
rect 1104 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8894 7642
rect 8946 7590 8958 7642
rect 9010 7590 9022 7642
rect 9074 7590 9086 7642
rect 9138 7590 12972 7642
rect 1104 7568 12972 7590
rect 1489 7531 1547 7537
rect 1489 7497 1501 7531
rect 1535 7528 1547 7531
rect 6454 7528 6460 7540
rect 1535 7500 6460 7528
rect 1535 7497 1547 7500
rect 1489 7491 1547 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 7650 7528 7656 7540
rect 6656 7500 7656 7528
rect 6656 7460 6684 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 2240 7432 6684 7460
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7392 1639 7395
rect 2130 7392 2136 7404
rect 1627 7364 2136 7392
rect 1627 7361 1639 7364
rect 1581 7355 1639 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2240 7401 2268 7432
rect 7282 7420 7288 7472
rect 7340 7460 7346 7472
rect 7469 7463 7527 7469
rect 7469 7460 7481 7463
rect 7340 7432 7481 7460
rect 7340 7420 7346 7432
rect 7469 7429 7481 7432
rect 7515 7460 7527 7463
rect 7515 7432 7788 7460
rect 7515 7429 7527 7432
rect 7469 7423 7527 7429
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 3145 7395 3203 7401
rect 3145 7392 3157 7395
rect 2556 7364 3157 7392
rect 2556 7352 2562 7364
rect 3145 7361 3157 7364
rect 3191 7361 3203 7395
rect 3145 7355 3203 7361
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3418 7392 3424 7404
rect 3292 7364 3424 7392
rect 3292 7352 3298 7364
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 7760 7401 7788 7432
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 11422 7392 11428 7404
rect 8619 7364 11428 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 2774 7324 2780 7336
rect 2740 7296 2780 7324
rect 2740 7284 2746 7296
rect 2774 7284 2780 7296
rect 2832 7324 2838 7336
rect 2869 7327 2927 7333
rect 2869 7324 2881 7327
rect 2832 7296 2881 7324
rect 2832 7284 2838 7296
rect 2869 7293 2881 7296
rect 2915 7293 2927 7327
rect 2869 7287 2927 7293
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 7926 7324 7932 7336
rect 7423 7296 7932 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 8018 7284 8024 7336
rect 8076 7324 8082 7336
rect 8294 7324 8300 7336
rect 8076 7296 8300 7324
rect 8076 7284 8082 7296
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 7466 7256 7472 7268
rect 3804 7228 7472 7256
rect 2133 7191 2191 7197
rect 2133 7157 2145 7191
rect 2179 7188 2191 7191
rect 3804 7188 3832 7228
rect 7466 7216 7472 7228
rect 7524 7216 7530 7268
rect 7653 7259 7711 7265
rect 7653 7225 7665 7259
rect 7699 7256 7711 7259
rect 9582 7256 9588 7268
rect 7699 7228 9588 7256
rect 7699 7225 7711 7228
rect 7653 7219 7711 7225
rect 9582 7216 9588 7228
rect 9640 7216 9646 7268
rect 2179 7160 3832 7188
rect 3881 7191 3939 7197
rect 2179 7157 2191 7160
rect 2133 7151 2191 7157
rect 3881 7157 3893 7191
rect 3927 7188 3939 7191
rect 8018 7188 8024 7200
rect 3927 7160 8024 7188
rect 3927 7157 3939 7160
rect 3881 7151 3939 7157
rect 8018 7148 8024 7160
rect 8076 7148 8082 7200
rect 8478 7188 8484 7200
rect 8439 7160 8484 7188
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 1104 7098 12972 7120
rect 1104 7046 2960 7098
rect 3012 7046 3024 7098
rect 3076 7046 3088 7098
rect 3140 7046 3152 7098
rect 3204 7046 6916 7098
rect 6968 7046 6980 7098
rect 7032 7046 7044 7098
rect 7096 7046 7108 7098
rect 7160 7046 10872 7098
rect 10924 7046 10936 7098
rect 10988 7046 11000 7098
rect 11052 7046 11064 7098
rect 11116 7046 12972 7098
rect 1104 7024 12972 7046
rect 2130 6944 2136 6996
rect 2188 6984 2194 6996
rect 6730 6984 6736 6996
rect 2188 6956 6736 6984
rect 2188 6944 2194 6956
rect 6730 6944 6736 6956
rect 6788 6984 6794 6996
rect 7466 6984 7472 6996
rect 6788 6956 7052 6984
rect 6788 6944 6794 6956
rect 7024 6928 7052 6956
rect 7208 6956 7472 6984
rect 7208 6928 7236 6956
rect 7466 6944 7472 6956
rect 7524 6984 7530 6996
rect 7742 6984 7748 6996
rect 7524 6956 7748 6984
rect 7524 6944 7530 6956
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 3418 6876 3424 6928
rect 3476 6916 3482 6928
rect 6181 6919 6239 6925
rect 6181 6916 6193 6919
rect 3476 6888 6193 6916
rect 3476 6876 3482 6888
rect 6181 6885 6193 6888
rect 6227 6885 6239 6919
rect 6181 6879 6239 6885
rect 6362 6876 6368 6928
rect 6420 6916 6426 6928
rect 6420 6888 6500 6916
rect 6420 6876 6426 6888
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 5534 6848 5540 6860
rect 2924 6820 5540 6848
rect 2924 6808 2930 6820
rect 5534 6808 5540 6820
rect 5592 6848 5598 6860
rect 6270 6848 6276 6860
rect 5592 6820 6276 6848
rect 5592 6808 5598 6820
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 2222 6780 2228 6792
rect 2183 6752 2228 6780
rect 2222 6740 2228 6752
rect 2280 6740 2286 6792
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2682 6780 2688 6792
rect 2547 6752 2688 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2682 6740 2688 6752
rect 2740 6780 2746 6792
rect 2740 6740 2774 6780
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4522 6780 4528 6792
rect 4304 6752 4528 6780
rect 4304 6740 4310 6752
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 6362 6780 6368 6792
rect 6323 6752 6368 6780
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6472 6789 6500 6888
rect 7006 6876 7012 6928
rect 7064 6876 7070 6928
rect 7190 6876 7196 6928
rect 7248 6876 7254 6928
rect 7300 6888 7604 6916
rect 7300 6848 7328 6888
rect 7466 6848 7472 6860
rect 6748 6820 7328 6848
rect 7392 6820 7472 6848
rect 6748 6789 6776 6820
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 7190 6780 7196 6792
rect 7151 6752 7196 6780
rect 6733 6743 6791 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7392 6789 7420 6820
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7576 6848 7604 6888
rect 8386 6848 8392 6860
rect 7576 6820 8392 6848
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 9214 6848 9220 6860
rect 8496 6820 9220 6848
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 7650 6780 7656 6792
rect 7607 6752 7656 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 2746 6712 2774 6740
rect 6086 6712 6092 6724
rect 2746 6684 6092 6712
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 6549 6715 6607 6721
rect 6549 6712 6561 6715
rect 6196 6684 6561 6712
rect 1489 6647 1547 6653
rect 1489 6613 1501 6647
rect 1535 6644 1547 6647
rect 1578 6644 1584 6656
rect 1535 6616 1584 6644
rect 1535 6613 1547 6616
rect 1489 6607 1547 6613
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 3970 6644 3976 6656
rect 3660 6616 3976 6644
rect 3660 6604 3666 6616
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 6196 6644 6224 6684
rect 6549 6681 6561 6684
rect 6595 6712 6607 6715
rect 7098 6712 7104 6724
rect 6595 6684 7104 6712
rect 6595 6681 6607 6684
rect 6549 6675 6607 6681
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 7469 6715 7527 6721
rect 7469 6681 7481 6715
rect 7515 6712 7527 6715
rect 8496 6712 8524 6820
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 12158 6848 12164 6860
rect 9646 6820 12164 6848
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 9646 6780 9674 6820
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 8628 6752 9674 6780
rect 8628 6740 8634 6752
rect 7515 6684 8524 6712
rect 7515 6681 7527 6684
rect 7469 6675 7527 6681
rect 8846 6672 8852 6724
rect 8904 6712 8910 6724
rect 8904 6684 9674 6712
rect 8904 6672 8910 6684
rect 4212 6616 6224 6644
rect 7745 6647 7803 6653
rect 4212 6604 4218 6616
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 9490 6644 9496 6656
rect 7791 6616 9496 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9646 6644 9674 6684
rect 10134 6672 10140 6724
rect 10192 6712 10198 6724
rect 10778 6712 10784 6724
rect 10192 6684 10784 6712
rect 10192 6672 10198 6684
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 12066 6712 12072 6724
rect 12027 6684 12072 6712
rect 12066 6672 12072 6684
rect 12124 6672 12130 6724
rect 10226 6644 10232 6656
rect 9646 6616 10232 6644
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 12158 6644 12164 6656
rect 12119 6616 12164 6644
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 1104 6554 12972 6576
rect 1104 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8894 6554
rect 8946 6502 8958 6554
rect 9010 6502 9022 6554
rect 9074 6502 9086 6554
rect 9138 6502 12972 6554
rect 1104 6480 12972 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 2593 6443 2651 6449
rect 2593 6409 2605 6443
rect 2639 6440 2651 6443
rect 3326 6440 3332 6452
rect 2639 6412 3332 6440
rect 2639 6409 2651 6412
rect 2593 6403 2651 6409
rect 1596 6372 1624 6403
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 5350 6440 5356 6452
rect 4571 6412 5356 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 4540 6372 4568 6403
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 6362 6400 6368 6452
rect 6420 6440 6426 6452
rect 8202 6440 8208 6452
rect 6420 6412 8208 6440
rect 6420 6400 6426 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9858 6440 9864 6452
rect 9784 6412 9864 6440
rect 7190 6372 7196 6384
rect 1596 6344 4568 6372
rect 5000 6344 7196 6372
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2740 6276 2789 6304
rect 2740 6264 2746 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 2866 6264 2872 6316
rect 2924 6304 2930 6316
rect 3145 6307 3203 6313
rect 2924 6276 2969 6304
rect 2924 6264 2930 6276
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 4062 6304 4068 6316
rect 3191 6276 4068 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 5000 6313 5028 6344
rect 7190 6332 7196 6344
rect 7248 6332 7254 6384
rect 7469 6375 7527 6381
rect 7469 6341 7481 6375
rect 7515 6372 7527 6375
rect 9784 6372 9812 6412
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 11514 6440 11520 6452
rect 10284 6412 11192 6440
rect 11475 6412 11520 6440
rect 10284 6400 10290 6412
rect 7515 6344 9812 6372
rect 11164 6372 11192 6412
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 11701 6443 11759 6449
rect 11701 6409 11713 6443
rect 11747 6409 11759 6443
rect 11701 6403 11759 6409
rect 11716 6372 11744 6403
rect 11164 6344 12112 6372
rect 7515 6341 7527 6344
rect 7469 6335 7527 6341
rect 4522 6307 4580 6313
rect 4522 6273 4534 6307
rect 4568 6304 4580 6307
rect 4985 6307 5043 6313
rect 4568 6276 4844 6304
rect 4568 6273 4580 6276
rect 4522 6267 4580 6273
rect 4816 6236 4844 6276
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5000 6236 5028 6267
rect 6086 6264 6092 6316
rect 6144 6304 6150 6316
rect 6638 6304 6644 6316
rect 6144 6276 6644 6304
rect 6144 6264 6150 6276
rect 6638 6264 6644 6276
rect 6696 6264 6702 6316
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7064 6276 7389 6304
rect 7064 6264 7070 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7650 6304 7656 6316
rect 7607 6276 7656 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6304 7803 6307
rect 8294 6304 8300 6316
rect 7791 6276 8300 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 9214 6304 9220 6316
rect 9175 6276 9220 6304
rect 9214 6264 9220 6276
rect 9272 6264 9278 6316
rect 9582 6264 9588 6316
rect 9640 6304 9646 6316
rect 9640 6302 9720 6304
rect 9766 6302 9772 6316
rect 9640 6276 9772 6302
rect 9640 6264 9646 6276
rect 9692 6274 9772 6276
rect 9766 6264 9772 6274
rect 9824 6264 9830 6316
rect 10410 6304 10416 6316
rect 10371 6276 10416 6304
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 12084 6313 12112 6344
rect 11698 6307 11756 6313
rect 11698 6273 11710 6307
rect 11744 6273 11756 6307
rect 11698 6267 11756 6273
rect 12069 6307 12127 6313
rect 12069 6273 12081 6307
rect 12115 6273 12127 6307
rect 12069 6267 12127 6273
rect 4816 6208 5028 6236
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 10042 6236 10048 6248
rect 9456 6208 10048 6236
rect 9456 6196 9462 6208
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10689 6239 10747 6245
rect 10689 6205 10701 6239
rect 10735 6236 10747 6239
rect 11238 6236 11244 6248
rect 10735 6208 11244 6236
rect 10735 6205 10747 6208
rect 10689 6199 10747 6205
rect 11238 6196 11244 6208
rect 11296 6196 11302 6248
rect 11514 6196 11520 6248
rect 11572 6236 11578 6248
rect 11716 6236 11744 6267
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 11572 6208 12173 6236
rect 11572 6196 11578 6208
rect 12161 6205 12173 6208
rect 12207 6205 12219 6239
rect 12161 6199 12219 6205
rect 2774 6128 2780 6180
rect 2832 6168 2838 6180
rect 3053 6171 3111 6177
rect 3053 6168 3065 6171
rect 2832 6140 3065 6168
rect 2832 6128 2838 6140
rect 3053 6137 3065 6140
rect 3099 6137 3111 6171
rect 8754 6168 8760 6180
rect 3053 6131 3111 6137
rect 3160 6140 8760 6168
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 3160 6100 3188 6140
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9125 6171 9183 6177
rect 9125 6168 9137 6171
rect 9088 6140 9137 6168
rect 9088 6128 9094 6140
rect 9125 6137 9137 6140
rect 9171 6168 9183 6171
rect 9766 6168 9772 6180
rect 9171 6140 9772 6168
rect 9171 6137 9183 6140
rect 9125 6131 9183 6137
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 10778 6128 10784 6180
rect 10836 6128 10842 6180
rect 2740 6072 3188 6100
rect 2740 6060 2746 6072
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 4341 6103 4399 6109
rect 4341 6100 4353 6103
rect 3660 6072 4353 6100
rect 3660 6060 3666 6072
rect 4341 6069 4353 6072
rect 4387 6100 4399 6103
rect 4798 6100 4804 6112
rect 4387 6072 4804 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4798 6060 4804 6072
rect 4856 6060 4862 6112
rect 4893 6103 4951 6109
rect 4893 6069 4905 6103
rect 4939 6100 4951 6103
rect 5350 6100 5356 6112
rect 4939 6072 5356 6100
rect 4939 6069 4951 6072
rect 4893 6063 4951 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 6788 6072 7205 6100
rect 6788 6060 6794 6072
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 7193 6063 7251 6069
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 10796 6100 10824 6128
rect 9723 6072 10824 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 1104 6010 12972 6032
rect 1104 5958 2960 6010
rect 3012 5958 3024 6010
rect 3076 5958 3088 6010
rect 3140 5958 3152 6010
rect 3204 5958 6916 6010
rect 6968 5958 6980 6010
rect 7032 5958 7044 6010
rect 7096 5958 7108 6010
rect 7160 5958 10872 6010
rect 10924 5958 10936 6010
rect 10988 5958 11000 6010
rect 11052 5958 11064 6010
rect 11116 5958 12972 6010
rect 1104 5936 12972 5958
rect 7282 5896 7288 5908
rect 4724 5868 7288 5896
rect 4522 5760 4528 5772
rect 4483 5732 4528 5760
rect 4522 5720 4528 5732
rect 4580 5720 4586 5772
rect 4430 5692 4436 5704
rect 4391 5664 4436 5692
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4724 5701 4752 5868
rect 7282 5856 7288 5868
rect 7340 5856 7346 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 10410 5896 10416 5908
rect 7708 5868 10416 5896
rect 7708 5856 7714 5868
rect 10410 5856 10416 5868
rect 10468 5896 10474 5908
rect 11698 5896 11704 5908
rect 10468 5868 11704 5896
rect 10468 5856 10474 5868
rect 11698 5856 11704 5868
rect 11756 5856 11762 5908
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5828 5043 5831
rect 5718 5828 5724 5840
rect 5031 5800 5724 5828
rect 5031 5797 5043 5800
rect 4985 5791 5043 5797
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 7116 5800 10272 5828
rect 6457 5763 6515 5769
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6638 5760 6644 5772
rect 6503 5732 6644 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6638 5720 6644 5732
rect 6696 5760 6702 5772
rect 6822 5760 6828 5772
rect 6696 5732 6828 5760
rect 6696 5720 6702 5732
rect 6822 5720 6828 5732
rect 6880 5720 6886 5772
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 5902 5692 5908 5704
rect 4847 5664 5908 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6178 5692 6184 5704
rect 6139 5664 6184 5692
rect 6178 5652 6184 5664
rect 6236 5652 6242 5704
rect 7116 5701 7144 5800
rect 7208 5732 8892 5760
rect 7208 5701 7236 5732
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 7449 5695 7507 5701
rect 7449 5661 7461 5695
rect 7495 5692 7507 5695
rect 8864 5692 8892 5732
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9582 5760 9588 5772
rect 9180 5732 9588 5760
rect 9180 5720 9186 5732
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 10244 5760 10272 5800
rect 10244 5732 10364 5760
rect 10134 5692 10140 5704
rect 7495 5682 7512 5692
rect 7576 5682 7972 5692
rect 7495 5664 7972 5682
rect 8864 5664 10140 5692
rect 7495 5661 7604 5664
rect 7449 5655 7604 5661
rect 7484 5654 7604 5655
rect 7285 5627 7343 5633
rect 7285 5593 7297 5627
rect 7331 5624 7343 5627
rect 7650 5624 7656 5636
rect 7331 5596 7656 5624
rect 7331 5593 7343 5596
rect 7285 5587 7343 5593
rect 7650 5584 7656 5596
rect 7708 5584 7714 5636
rect 7944 5624 7972 5664
rect 10134 5652 10140 5664
rect 10192 5652 10198 5704
rect 10226 5624 10232 5636
rect 7944 5596 10232 5624
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 6917 5559 6975 5565
rect 6917 5556 6929 5559
rect 5592 5528 6929 5556
rect 5592 5516 5598 5528
rect 6917 5525 6929 5528
rect 6963 5525 6975 5559
rect 6917 5519 6975 5525
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 9861 5559 9919 5565
rect 9861 5556 9873 5559
rect 8352 5528 9873 5556
rect 8352 5516 8358 5528
rect 9861 5525 9873 5528
rect 9907 5525 9919 5559
rect 10336 5556 10364 5732
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12032 5732 12204 5760
rect 12032 5720 12038 5732
rect 10594 5652 10600 5704
rect 10652 5692 10658 5704
rect 10870 5692 10876 5704
rect 10652 5664 10697 5692
rect 10831 5664 10876 5692
rect 10652 5652 10658 5664
rect 10870 5652 10876 5664
rect 10928 5692 10934 5704
rect 11238 5692 11244 5704
rect 10928 5664 11244 5692
rect 10928 5652 10934 5664
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 12176 5701 12204 5732
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 10778 5584 10784 5636
rect 10836 5624 10842 5636
rect 11793 5627 11851 5633
rect 11793 5624 11805 5627
rect 10836 5596 11805 5624
rect 10836 5584 10842 5596
rect 11793 5593 11805 5596
rect 11839 5593 11851 5627
rect 11793 5587 11851 5593
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 12032 5596 12077 5624
rect 12032 5584 12038 5596
rect 12176 5556 12204 5655
rect 10336 5528 12204 5556
rect 9861 5519 9919 5525
rect 1104 5466 12972 5488
rect 1104 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8894 5466
rect 8946 5414 8958 5466
rect 9010 5414 9022 5466
rect 9074 5414 9086 5466
rect 9138 5414 12972 5466
rect 1104 5392 12972 5414
rect 3237 5355 3295 5361
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 5810 5352 5816 5364
rect 3283 5324 5816 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 5810 5312 5816 5324
rect 5868 5312 5874 5364
rect 5902 5312 5908 5364
rect 5960 5352 5966 5364
rect 7926 5352 7932 5364
rect 5960 5324 7932 5352
rect 5960 5312 5966 5324
rect 7926 5312 7932 5324
rect 7984 5352 7990 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 7984 5324 12265 5352
rect 7984 5312 7990 5324
rect 12253 5321 12265 5324
rect 12299 5321 12311 5355
rect 12253 5315 12311 5321
rect 5169 5287 5227 5293
rect 5169 5253 5181 5287
rect 5215 5284 5227 5287
rect 7466 5284 7472 5296
rect 5215 5256 7472 5284
rect 5215 5253 5227 5256
rect 5169 5247 5227 5253
rect 7466 5244 7472 5256
rect 7524 5244 7530 5296
rect 10594 5244 10600 5296
rect 10652 5284 10658 5296
rect 10870 5284 10876 5296
rect 10652 5256 10876 5284
rect 10652 5244 10658 5256
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11882 5284 11888 5296
rect 11843 5256 11888 5284
rect 11882 5244 11888 5256
rect 11940 5244 11946 5296
rect 3418 5216 3424 5228
rect 3379 5188 3424 5216
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 3510 5176 3516 5228
rect 3568 5216 3574 5228
rect 3789 5219 3847 5225
rect 3568 5188 3613 5216
rect 3568 5176 3574 5188
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 4154 5216 4160 5228
rect 3835 5188 4160 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5810 5216 5816 5228
rect 5307 5188 5816 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 6604 5188 6649 5216
rect 6604 5176 6610 5188
rect 7834 5176 7840 5228
rect 7892 5216 7898 5228
rect 11238 5216 11244 5228
rect 7892 5188 11244 5216
rect 7892 5176 7898 5188
rect 11238 5176 11244 5188
rect 11296 5176 11302 5228
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11563 5188 11713 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12069 5179 12127 5185
rect 3697 5151 3755 5157
rect 3697 5117 3709 5151
rect 3743 5148 3755 5151
rect 5902 5148 5908 5160
rect 3743 5120 5908 5148
rect 3743 5117 3755 5120
rect 3697 5111 3755 5117
rect 5902 5108 5908 5120
rect 5960 5108 5966 5160
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 11992 5148 12020 5179
rect 9272 5120 12020 5148
rect 9272 5108 9278 5120
rect 6457 5083 6515 5089
rect 6457 5049 6469 5083
rect 6503 5080 6515 5083
rect 10318 5080 10324 5092
rect 6503 5052 10324 5080
rect 6503 5049 6515 5052
rect 6457 5043 6515 5049
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 11974 5080 11980 5092
rect 11296 5052 11980 5080
rect 11296 5040 11302 5052
rect 11974 5040 11980 5052
rect 12032 5080 12038 5092
rect 12084 5080 12112 5179
rect 12032 5052 12112 5080
rect 12032 5040 12038 5052
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 4580 4984 11529 5012
rect 4580 4972 4586 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 1104 4922 12972 4944
rect 1104 4870 2960 4922
rect 3012 4870 3024 4922
rect 3076 4870 3088 4922
rect 3140 4870 3152 4922
rect 3204 4870 6916 4922
rect 6968 4870 6980 4922
rect 7032 4870 7044 4922
rect 7096 4870 7108 4922
rect 7160 4870 10872 4922
rect 10924 4870 10936 4922
rect 10988 4870 11000 4922
rect 11052 4870 11064 4922
rect 11116 4870 12972 4922
rect 1104 4848 12972 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2222 4808 2228 4820
rect 2087 4780 2228 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4985 4811 5043 4817
rect 4985 4808 4997 4811
rect 4672 4780 4997 4808
rect 4672 4768 4678 4780
rect 4985 4777 4997 4780
rect 5031 4777 5043 4811
rect 5534 4808 5540 4820
rect 4985 4771 5043 4777
rect 5092 4780 5540 4808
rect 2593 4743 2651 4749
rect 2593 4740 2605 4743
rect 2148 4712 2605 4740
rect 2148 4468 2176 4712
rect 2593 4709 2605 4712
rect 2639 4740 2651 4743
rect 5092 4740 5120 4780
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 8386 4808 8392 4820
rect 5960 4780 8392 4808
rect 5960 4768 5966 4780
rect 8386 4768 8392 4780
rect 8444 4808 8450 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 8444 4780 9413 4808
rect 8444 4768 8450 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 2639 4712 5120 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 5994 4700 6000 4752
rect 6052 4740 6058 4752
rect 11241 4743 11299 4749
rect 11241 4740 11253 4743
rect 6052 4712 11253 4740
rect 6052 4700 6058 4712
rect 11241 4709 11253 4712
rect 11287 4709 11299 4743
rect 11241 4703 11299 4709
rect 2685 4675 2743 4681
rect 2685 4672 2697 4675
rect 2237 4644 2697 4672
rect 2237 4613 2265 4644
rect 2685 4641 2697 4644
rect 2731 4672 2743 4675
rect 3602 4672 3608 4684
rect 2731 4644 3608 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 3602 4632 3608 4644
rect 3660 4632 3666 4684
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 8536 4644 11836 4672
rect 8536 4632 8542 4644
rect 2222 4607 2280 4613
rect 2222 4573 2234 4607
rect 2268 4573 2280 4607
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 2222 4567 2280 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 3878 4564 3884 4616
rect 3936 4604 3942 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3936 4576 3985 4604
rect 3936 4564 3942 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4061 4607 4119 4613
rect 4061 4573 4073 4607
rect 4107 4573 4119 4607
rect 4061 4567 4119 4573
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4246 4604 4252 4616
rect 4203 4576 4252 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 2225 4471 2283 4477
rect 2225 4468 2237 4471
rect 2148 4440 2237 4468
rect 2225 4437 2237 4440
rect 2271 4437 2283 4471
rect 2225 4431 2283 4437
rect 3970 4428 3976 4480
rect 4028 4468 4034 4480
rect 4080 4468 4108 4567
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5997 4607 6055 4613
rect 5997 4573 6009 4607
rect 6043 4604 6055 4607
rect 6638 4604 6644 4616
rect 6043 4576 6644 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 5736 4536 5764 4567
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 8260 4576 9505 4604
rect 8260 4564 8266 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 11422 4604 11428 4616
rect 11383 4576 11428 4604
rect 9493 4567 9551 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11808 4613 11836 4644
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 7282 4536 7288 4548
rect 5736 4508 7288 4536
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 11514 4536 11520 4548
rect 11475 4508 11520 4536
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 4028 4440 4108 4468
rect 4341 4471 4399 4477
rect 4028 4428 4034 4440
rect 4341 4437 4353 4471
rect 4387 4468 4399 4471
rect 5258 4468 5264 4480
rect 4387 4440 5264 4468
rect 4387 4437 4399 4440
rect 4341 4431 4399 4437
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 11882 4468 11888 4480
rect 8444 4440 11888 4468
rect 8444 4428 8450 4440
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 1104 4378 12972 4400
rect 1104 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8894 4378
rect 8946 4326 8958 4378
rect 9010 4326 9022 4378
rect 9074 4326 9086 4378
rect 9138 4326 12972 4378
rect 1104 4304 12972 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3973 4267 4031 4273
rect 3973 4264 3985 4267
rect 2832 4236 3985 4264
rect 2832 4224 2838 4236
rect 3973 4233 3985 4236
rect 4019 4233 4031 4267
rect 3973 4227 4031 4233
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 8386 4264 8392 4276
rect 4764 4236 8392 4264
rect 4764 4224 4770 4236
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 8662 4224 8668 4276
rect 8720 4264 8726 4276
rect 8941 4267 8999 4273
rect 8941 4264 8953 4267
rect 8720 4236 8953 4264
rect 8720 4224 8726 4236
rect 8941 4233 8953 4236
rect 8987 4264 8999 4267
rect 8987 4236 11744 4264
rect 8987 4233 8999 4236
rect 8941 4227 8999 4233
rect 1949 4199 2007 4205
rect 1949 4165 1961 4199
rect 1995 4196 2007 4199
rect 8294 4196 8300 4208
rect 1995 4168 8300 4196
rect 1995 4165 2007 4168
rect 1949 4159 2007 4165
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 8404 4196 8432 4224
rect 11716 4205 11744 4236
rect 11701 4199 11759 4205
rect 8404 4168 8708 4196
rect 4065 4131 4123 4137
rect 4065 4097 4077 4131
rect 4111 4128 4123 4131
rect 5350 4128 5356 4140
rect 4111 4100 5356 4128
rect 4111 4097 4123 4100
rect 4065 4091 4123 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 8680 4128 8708 4168
rect 10060 4168 10916 4196
rect 8944 4131 9002 4137
rect 8944 4128 8956 4131
rect 7800 4100 8616 4128
rect 8680 4100 8956 4128
rect 7800 4088 7806 4100
rect 8386 4020 8392 4072
rect 8444 4060 8450 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8444 4032 8493 4060
rect 8444 4020 8450 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 8588 4060 8616 4100
rect 8944 4097 8956 4100
rect 8990 4097 9002 4131
rect 10060 4128 10088 4168
rect 8944 4091 9002 4097
rect 9140 4100 10088 4128
rect 10137 4131 10195 4137
rect 9140 4060 9168 4100
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10318 4128 10324 4140
rect 10183 4100 10324 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10560 4100 10824 4128
rect 10560 4088 10566 4100
rect 8588 4032 9168 4060
rect 8481 4023 8539 4029
rect 9490 4020 9496 4072
rect 9548 4060 9554 4072
rect 10796 4069 10824 4100
rect 10888 4069 10916 4168
rect 11701 4165 11713 4199
rect 11747 4165 11759 4199
rect 11882 4196 11888 4208
rect 11843 4168 11888 4196
rect 11701 4159 11759 4165
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 9548 4032 10609 4060
rect 9548 4020 9554 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10781 4063 10839 4069
rect 10781 4029 10793 4063
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 10873 4063 10931 4069
rect 10873 4029 10885 4063
rect 10919 4029 10931 4063
rect 10873 4023 10931 4029
rect 7466 3952 7472 4004
rect 7524 3992 7530 4004
rect 9125 3995 9183 4001
rect 7524 3964 8708 3992
rect 7524 3952 7530 3964
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 8570 3924 8576 3936
rect 8531 3896 8576 3924
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8680 3924 8708 3964
rect 9125 3961 9137 3995
rect 9171 3992 9183 3995
rect 9398 3992 9404 4004
rect 9171 3964 9404 3992
rect 9171 3961 9183 3964
rect 9125 3955 9183 3961
rect 9398 3952 9404 3964
rect 9456 3952 9462 4004
rect 9950 3992 9956 4004
rect 9911 3964 9956 3992
rect 9950 3952 9956 3964
rect 10008 3952 10014 4004
rect 10980 3992 11008 4091
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 12069 4063 12127 4069
rect 12069 4060 12081 4063
rect 11848 4032 12081 4060
rect 11848 4020 11854 4032
rect 12069 4029 12081 4032
rect 12115 4029 12127 4063
rect 12069 4023 12127 4029
rect 10060 3964 11008 3992
rect 10060 3924 10088 3964
rect 8680 3896 10088 3924
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 10781 3927 10839 3933
rect 10781 3924 10793 3927
rect 10744 3896 10793 3924
rect 10744 3884 10750 3896
rect 10781 3893 10793 3896
rect 10827 3893 10839 3927
rect 10781 3887 10839 3893
rect 1104 3834 12972 3856
rect 1104 3782 2960 3834
rect 3012 3782 3024 3834
rect 3076 3782 3088 3834
rect 3140 3782 3152 3834
rect 3204 3782 6916 3834
rect 6968 3782 6980 3834
rect 7032 3782 7044 3834
rect 7096 3782 7108 3834
rect 7160 3782 10872 3834
rect 10924 3782 10936 3834
rect 10988 3782 11000 3834
rect 11052 3782 11064 3834
rect 11116 3782 12972 3834
rect 1104 3760 12972 3782
rect 5626 3680 5632 3732
rect 5684 3720 5690 3732
rect 7009 3723 7067 3729
rect 7009 3720 7021 3723
rect 5684 3692 7021 3720
rect 5684 3680 5690 3692
rect 7009 3689 7021 3692
rect 7055 3689 7067 3723
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 7009 3683 7067 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10410 3680 10416 3732
rect 10468 3720 10474 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10468 3692 10701 3720
rect 10468 3680 10474 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 1581 3655 1639 3661
rect 1581 3621 1593 3655
rect 1627 3652 1639 3655
rect 6454 3652 6460 3664
rect 1627 3624 6460 3652
rect 1627 3621 1639 3624
rect 1581 3615 1639 3621
rect 6454 3612 6460 3624
rect 6512 3612 6518 3664
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 6779 3556 7297 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 7285 3553 7297 3556
rect 7331 3584 7343 3587
rect 9306 3584 9312 3596
rect 7331 3556 9312 3584
rect 7331 3553 7343 3556
rect 7285 3547 7343 3553
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 9548 3556 9597 3584
rect 9548 3544 9554 3556
rect 9585 3553 9597 3556
rect 9631 3584 9643 3587
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9631 3556 10149 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 11974 3584 11980 3596
rect 11935 3556 11980 3584
rect 10137 3547 10195 3553
rect 11974 3544 11980 3556
rect 12032 3544 12038 3596
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 6840 3488 7113 3516
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6840 3457 6868 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 9953 3519 10011 3525
rect 9953 3485 9965 3519
rect 9999 3485 10011 3519
rect 9953 3479 10011 3485
rect 6825 3451 6883 3457
rect 6825 3448 6837 3451
rect 5776 3420 6837 3448
rect 5776 3408 5782 3420
rect 6825 3417 6837 3420
rect 6871 3417 6883 3451
rect 6825 3411 6883 3417
rect 9677 3451 9735 3457
rect 9677 3417 9689 3451
rect 9723 3448 9735 3451
rect 9968 3448 9996 3479
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10100 3488 10609 3516
rect 10100 3476 10106 3488
rect 10597 3485 10609 3488
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 12253 3519 12311 3525
rect 12253 3485 12265 3519
rect 12299 3516 12311 3519
rect 12894 3516 12900 3528
rect 12299 3488 12900 3516
rect 12299 3485 12311 3488
rect 12253 3479 12311 3485
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 10502 3448 10508 3460
rect 9723 3420 10508 3448
rect 9723 3417 9735 3420
rect 9677 3411 9735 3417
rect 10502 3408 10508 3420
rect 10560 3408 10566 3460
rect 1104 3290 12972 3312
rect 1104 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8894 3290
rect 8946 3238 8958 3290
rect 9010 3238 9022 3290
rect 9074 3238 9086 3290
rect 9138 3238 12972 3290
rect 1104 3216 12972 3238
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 8573 3179 8631 3185
rect 8573 3176 8585 3179
rect 7340 3148 8585 3176
rect 7340 3136 7346 3148
rect 8573 3145 8585 3148
rect 8619 3145 8631 3179
rect 8573 3139 8631 3145
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 12158 3176 12164 3188
rect 9732 3148 9777 3176
rect 12119 3148 12164 3176
rect 9732 3136 9738 3148
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 6270 3068 6276 3120
rect 6328 3108 6334 3120
rect 8481 3111 8539 3117
rect 8481 3108 8493 3111
rect 6328 3080 8493 3108
rect 6328 3068 6334 3080
rect 8481 3077 8493 3080
rect 8527 3077 8539 3111
rect 8481 3071 8539 3077
rect 14 3000 20 3052
rect 72 3040 78 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 72 3012 1409 3040
rect 72 3000 78 3012
rect 1397 3009 1409 3012
rect 1443 3009 1455 3043
rect 8496 3040 8524 3071
rect 10594 3068 10600 3120
rect 10652 3108 10658 3120
rect 10652 3080 10732 3108
rect 10652 3068 10658 3080
rect 8757 3043 8815 3049
rect 8757 3040 8769 3043
rect 8496 3012 8769 3040
rect 1397 3003 1455 3009
rect 8757 3009 8769 3012
rect 8803 3009 8815 3043
rect 8757 3003 8815 3009
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 10704 3049 10732 3080
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 12069 3111 12127 3117
rect 12069 3108 12081 3111
rect 11388 3080 12081 3108
rect 11388 3068 11394 3080
rect 12069 3077 12081 3080
rect 12115 3077 12127 3111
rect 12069 3071 12127 3077
rect 8941 3043 8999 3049
rect 8941 3040 8953 3043
rect 8904 3012 8953 3040
rect 8904 3000 8910 3012
rect 8941 3009 8953 3012
rect 8987 3009 8999 3043
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 8941 3003 8999 3009
rect 9324 3012 10425 3040
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 8864 2972 8892 3000
rect 8435 2944 8892 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 9214 2904 9220 2916
rect 1627 2876 9220 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 3694 2796 3700 2848
rect 3752 2836 3758 2848
rect 9324 2836 9352 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 3752 2808 9352 2836
rect 3752 2796 3758 2808
rect 1104 2746 12972 2768
rect 1104 2694 2960 2746
rect 3012 2694 3024 2746
rect 3076 2694 3088 2746
rect 3140 2694 3152 2746
rect 3204 2694 6916 2746
rect 6968 2694 6980 2746
rect 7032 2694 7044 2746
rect 7096 2694 7108 2746
rect 7160 2694 10872 2746
rect 10924 2694 10936 2746
rect 10988 2694 11000 2746
rect 11052 2694 11064 2746
rect 11116 2694 12972 2746
rect 1104 2672 12972 2694
rect 4157 2635 4215 2641
rect 4157 2601 4169 2635
rect 4203 2632 4215 2635
rect 10781 2635 10839 2641
rect 4203 2604 10732 2632
rect 4203 2601 4215 2604
rect 4157 2595 4215 2601
rect 3789 2567 3847 2573
rect 3789 2533 3801 2567
rect 3835 2564 3847 2567
rect 3835 2536 5672 2564
rect 3835 2533 3847 2536
rect 3789 2527 3847 2533
rect 5644 2496 5672 2536
rect 6546 2524 6552 2576
rect 6604 2564 6610 2576
rect 6733 2567 6791 2573
rect 6733 2564 6745 2567
rect 6604 2536 6745 2564
rect 6604 2524 6610 2536
rect 6733 2533 6745 2536
rect 6779 2533 6791 2567
rect 7374 2564 7380 2576
rect 6733 2527 6791 2533
rect 6886 2536 7380 2564
rect 6886 2496 6914 2536
rect 7374 2524 7380 2536
rect 7432 2524 7438 2576
rect 8570 2524 8576 2576
rect 8628 2564 8634 2576
rect 9309 2567 9367 2573
rect 9309 2564 9321 2567
rect 8628 2536 9321 2564
rect 8628 2524 8634 2536
rect 9309 2533 9321 2536
rect 9355 2533 9367 2567
rect 9309 2527 9367 2533
rect 9674 2496 9680 2508
rect 1964 2468 5580 2496
rect 5644 2468 6914 2496
rect 7392 2468 9680 2496
rect 1964 2437 1992 2468
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2397 2007 2431
rect 1949 2391 2007 2397
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2428 2927 2431
rect 3789 2431 3847 2437
rect 3789 2428 3801 2431
rect 2915 2400 3801 2428
rect 2915 2397 2927 2400
rect 2869 2391 2927 2397
rect 3789 2397 3801 2400
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 5442 2428 5448 2440
rect 5403 2400 5448 2428
rect 3973 2391 4031 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1765 2363 1823 2369
rect 1765 2360 1777 2363
rect 1360 2332 1777 2360
rect 1360 2320 1366 2332
rect 1765 2329 1777 2332
rect 1811 2329 1823 2363
rect 1765 2323 1823 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 2685 2363 2743 2369
rect 2685 2360 2697 2363
rect 2648 2332 2697 2360
rect 2648 2320 2654 2332
rect 2685 2329 2697 2332
rect 2731 2329 2743 2363
rect 5258 2360 5264 2372
rect 5219 2332 5264 2360
rect 2685 2323 2743 2329
rect 5258 2320 5264 2332
rect 5316 2320 5322 2372
rect 5552 2360 5580 2468
rect 6454 2388 6460 2440
rect 6512 2428 6518 2440
rect 7392 2437 7420 2468
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 10704 2496 10732 2604
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 11422 2632 11428 2644
rect 10827 2604 11428 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 11606 2592 11612 2644
rect 11664 2632 11670 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11664 2604 11713 2632
rect 11664 2592 11670 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 11514 2524 11520 2576
rect 11572 2524 11578 2576
rect 11532 2496 11560 2524
rect 10704 2468 11652 2496
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6512 2400 6561 2428
rect 6512 2388 6518 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 8018 2428 8024 2440
rect 7979 2400 8024 2428
rect 7377 2391 7435 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 9125 2431 9183 2437
rect 9125 2397 9137 2431
rect 9171 2428 9183 2431
rect 9214 2428 9220 2440
rect 9171 2400 9220 2428
rect 9171 2397 9183 2400
rect 9125 2391 9183 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10410 2428 10416 2440
rect 10367 2400 10416 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2428 11023 2431
rect 11514 2428 11520 2440
rect 11011 2400 11520 2428
rect 11011 2397 11023 2400
rect 10965 2391 11023 2397
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 11624 2437 11652 2468
rect 11609 2431 11667 2437
rect 11609 2397 11621 2431
rect 11655 2397 11667 2431
rect 11609 2391 11667 2397
rect 5552 2332 7604 2360
rect 7193 2295 7251 2301
rect 7193 2261 7205 2295
rect 7239 2292 7251 2295
rect 7466 2292 7472 2304
rect 7239 2264 7472 2292
rect 7239 2261 7251 2264
rect 7193 2255 7251 2261
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 7576 2292 7604 2332
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 7837 2363 7895 2369
rect 7837 2360 7849 2363
rect 7800 2332 7849 2360
rect 7800 2320 7806 2332
rect 7837 2329 7849 2332
rect 7883 2329 7895 2363
rect 7837 2323 7895 2329
rect 8110 2292 8116 2304
rect 7576 2264 8116 2292
rect 8110 2252 8116 2264
rect 8168 2252 8174 2304
rect 10134 2292 10140 2304
rect 10095 2264 10140 2292
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 1104 2202 12972 2224
rect 1104 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8894 2202
rect 8946 2150 8958 2202
rect 9010 2150 9022 2202
rect 9074 2150 9086 2202
rect 9138 2150 12972 2202
rect 1104 2128 12972 2150
rect 9582 2048 9588 2100
rect 9640 2088 9646 2100
rect 10134 2088 10140 2100
rect 9640 2060 10140 2088
rect 9640 2048 9646 2060
rect 10134 2048 10140 2060
rect 10192 2048 10198 2100
<< via1 >>
rect 8024 13676 8076 13728
rect 9772 13676 9824 13728
rect 2960 13574 3012 13626
rect 3024 13574 3076 13626
rect 3088 13574 3140 13626
rect 3152 13574 3204 13626
rect 6916 13574 6968 13626
rect 6980 13574 7032 13626
rect 7044 13574 7096 13626
rect 7108 13574 7160 13626
rect 10872 13574 10924 13626
rect 10936 13574 10988 13626
rect 11000 13574 11052 13626
rect 11064 13574 11116 13626
rect 5356 13472 5408 13524
rect 3424 13404 3476 13456
rect 1768 13379 1820 13388
rect 1768 13345 1777 13379
rect 1777 13345 1811 13379
rect 1811 13345 1820 13379
rect 1768 13336 1820 13345
rect 1860 13336 1912 13388
rect 2780 13268 2832 13320
rect 4436 13268 4488 13320
rect 5724 13404 5776 13456
rect 7288 13404 7340 13456
rect 1492 13200 1544 13252
rect 5448 13200 5500 13252
rect 8300 13268 8352 13320
rect 10968 13379 11020 13388
rect 9772 13268 9824 13320
rect 10968 13345 10977 13379
rect 10977 13345 11011 13379
rect 11011 13345 11020 13379
rect 10968 13336 11020 13345
rect 11888 13311 11940 13320
rect 9588 13200 9640 13252
rect 11888 13277 11897 13311
rect 11897 13277 11931 13311
rect 11931 13277 11940 13311
rect 11888 13268 11940 13277
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 12072 13200 12124 13252
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 4528 13132 4580 13184
rect 5264 13132 5316 13184
rect 6552 13132 6604 13184
rect 7472 13132 7524 13184
rect 8300 13132 8352 13184
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 8894 13030 8946 13082
rect 8958 13030 9010 13082
rect 9022 13030 9074 13082
rect 9086 13030 9138 13082
rect 2688 12928 2740 12980
rect 9864 12928 9916 12980
rect 11796 12928 11848 12980
rect 11980 12928 12032 12980
rect 572 12860 624 12912
rect 3424 12835 3476 12844
rect 3424 12801 3433 12835
rect 3433 12801 3467 12835
rect 3467 12801 3476 12835
rect 3424 12792 3476 12801
rect 3976 12903 4028 12912
rect 3976 12869 3985 12903
rect 3985 12869 4019 12903
rect 4019 12869 4028 12903
rect 3976 12860 4028 12869
rect 4620 12860 4672 12912
rect 5540 12860 5592 12912
rect 4344 12792 4396 12844
rect 4712 12792 4764 12844
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 8300 12792 8352 12844
rect 9956 12860 10008 12912
rect 12164 12860 12216 12912
rect 9312 12835 9364 12844
rect 9312 12801 9321 12835
rect 9321 12801 9355 12835
rect 9355 12801 9364 12835
rect 9312 12792 9364 12801
rect 9772 12792 9824 12844
rect 11704 12835 11756 12844
rect 11704 12801 11710 12835
rect 11710 12801 11744 12835
rect 11744 12801 11756 12835
rect 11704 12792 11756 12801
rect 11888 12792 11940 12844
rect 4252 12656 4304 12708
rect 7288 12656 7340 12708
rect 7564 12699 7616 12708
rect 7564 12665 7573 12699
rect 7573 12665 7607 12699
rect 7607 12665 7616 12699
rect 7564 12656 7616 12665
rect 10324 12656 10376 12708
rect 10416 12656 10468 12708
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 4160 12588 4212 12597
rect 10508 12588 10560 12640
rect 11980 12588 12032 12640
rect 2960 12486 3012 12538
rect 3024 12486 3076 12538
rect 3088 12486 3140 12538
rect 3152 12486 3204 12538
rect 6916 12486 6968 12538
rect 6980 12486 7032 12538
rect 7044 12486 7096 12538
rect 7108 12486 7160 12538
rect 10872 12486 10924 12538
rect 10936 12486 10988 12538
rect 11000 12486 11052 12538
rect 11064 12486 11116 12538
rect 3884 12384 3936 12436
rect 3700 12316 3752 12368
rect 10600 12384 10652 12436
rect 10784 12316 10836 12368
rect 4160 12248 4212 12300
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 1768 12112 1820 12164
rect 2412 12087 2464 12096
rect 2412 12053 2421 12087
rect 2421 12053 2455 12087
rect 2455 12053 2464 12087
rect 2412 12044 2464 12053
rect 4068 12180 4120 12232
rect 8392 12248 8444 12300
rect 9496 12248 9548 12300
rect 13452 12248 13504 12300
rect 4344 12223 4396 12232
rect 4344 12189 4353 12223
rect 4353 12189 4387 12223
rect 4387 12189 4396 12223
rect 4344 12180 4396 12189
rect 6000 12180 6052 12232
rect 9220 12180 9272 12232
rect 4436 12112 4488 12164
rect 5816 12044 5868 12096
rect 7656 12044 7708 12096
rect 10048 12112 10100 12164
rect 12072 12044 12124 12096
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 8894 11942 8946 11994
rect 8958 11942 9010 11994
rect 9022 11942 9074 11994
rect 9086 11942 9138 11994
rect 9312 11840 9364 11892
rect 9680 11772 9732 11824
rect 1400 11679 1452 11688
rect 1400 11645 1409 11679
rect 1409 11645 1443 11679
rect 1443 11645 1452 11679
rect 1400 11636 1452 11645
rect 6368 11704 6420 11756
rect 6920 11747 6972 11756
rect 5724 11636 5776 11688
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 8300 11704 8352 11756
rect 8392 11704 8444 11756
rect 10692 11704 10744 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 11704 11747 11756 11756
rect 10784 11704 10836 11713
rect 11704 11713 11713 11747
rect 11713 11713 11747 11747
rect 11747 11713 11756 11747
rect 11704 11704 11756 11713
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 8024 11636 8076 11688
rect 6460 11568 6512 11620
rect 3608 11500 3660 11552
rect 3884 11500 3936 11552
rect 3976 11500 4028 11552
rect 6736 11500 6788 11552
rect 9220 11500 9272 11552
rect 9772 11500 9824 11552
rect 2960 11398 3012 11450
rect 3024 11398 3076 11450
rect 3088 11398 3140 11450
rect 3152 11398 3204 11450
rect 6916 11398 6968 11450
rect 6980 11398 7032 11450
rect 7044 11398 7096 11450
rect 7108 11398 7160 11450
rect 10872 11398 10924 11450
rect 10936 11398 10988 11450
rect 11000 11398 11052 11450
rect 11064 11398 11116 11450
rect 4712 11339 4764 11348
rect 4712 11305 4721 11339
rect 4721 11305 4755 11339
rect 4755 11305 4764 11339
rect 4712 11296 4764 11305
rect 9772 11296 9824 11348
rect 10232 11296 10284 11348
rect 3884 11228 3936 11280
rect 4712 11160 4764 11212
rect 5264 11160 5316 11212
rect 3424 11092 3476 11144
rect 4068 11092 4120 11144
rect 9220 11228 9272 11280
rect 9312 11228 9364 11280
rect 3792 11024 3844 11076
rect 7564 11160 7616 11212
rect 11152 11160 11204 11212
rect 6460 11092 6512 11144
rect 10600 11092 10652 11144
rect 12256 11135 12308 11144
rect 5264 10956 5316 11008
rect 7288 11024 7340 11076
rect 8208 11024 8260 11076
rect 10232 11024 10284 11076
rect 11152 11067 11204 11076
rect 11152 11033 11161 11067
rect 11161 11033 11195 11067
rect 11195 11033 11204 11067
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 11152 11024 11204 11033
rect 10416 10956 10468 11008
rect 10692 10956 10744 11008
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 8894 10854 8946 10906
rect 8958 10854 9010 10906
rect 9022 10854 9074 10906
rect 9086 10854 9138 10906
rect 5540 10752 5592 10804
rect 6368 10752 6420 10804
rect 9404 10752 9456 10804
rect 4712 10684 4764 10736
rect 7748 10684 7800 10736
rect 11796 10616 11848 10668
rect 8668 10548 8720 10600
rect 6184 10480 6236 10532
rect 6276 10480 6328 10532
rect 11888 10480 11940 10532
rect 7380 10412 7432 10464
rect 7564 10412 7616 10464
rect 2960 10310 3012 10362
rect 3024 10310 3076 10362
rect 3088 10310 3140 10362
rect 3152 10310 3204 10362
rect 6916 10310 6968 10362
rect 6980 10310 7032 10362
rect 7044 10310 7096 10362
rect 7108 10310 7160 10362
rect 10872 10310 10924 10362
rect 10936 10310 10988 10362
rect 11000 10310 11052 10362
rect 11064 10310 11116 10362
rect 3792 10208 3844 10260
rect 4344 10208 4396 10260
rect 7472 10208 7524 10260
rect 9956 10208 10008 10260
rect 12164 10208 12216 10260
rect 3332 10140 3384 10192
rect 4344 10004 4396 10056
rect 4528 10047 4580 10056
rect 4528 10013 4537 10047
rect 4537 10013 4571 10047
rect 4571 10013 4580 10047
rect 9496 10140 9548 10192
rect 4528 10004 4580 10013
rect 9864 10004 9916 10056
rect 10968 10047 11020 10056
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 4068 9868 4120 9920
rect 5540 9868 5592 9920
rect 8760 9868 8812 9920
rect 10232 9868 10284 9920
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 8894 9766 8946 9818
rect 8958 9766 9010 9818
rect 9022 9766 9074 9818
rect 9086 9766 9138 9818
rect 1952 9664 2004 9716
rect 6276 9664 6328 9716
rect 6368 9664 6420 9716
rect 10968 9664 11020 9716
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 11520 9596 11572 9648
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10048 9435 10100 9444
rect 6736 9367 6788 9376
rect 6736 9333 6745 9367
rect 6745 9333 6779 9367
rect 6779 9333 6788 9367
rect 6736 9324 6788 9333
rect 7380 9324 7432 9376
rect 10048 9401 10057 9435
rect 10057 9401 10091 9435
rect 10091 9401 10100 9435
rect 10048 9392 10100 9401
rect 9312 9324 9364 9376
rect 10692 9324 10744 9376
rect 11244 9324 11296 9376
rect 2960 9222 3012 9274
rect 3024 9222 3076 9274
rect 3088 9222 3140 9274
rect 3152 9222 3204 9274
rect 6916 9222 6968 9274
rect 6980 9222 7032 9274
rect 7044 9222 7096 9274
rect 7108 9222 7160 9274
rect 10872 9222 10924 9274
rect 10936 9222 10988 9274
rect 11000 9222 11052 9274
rect 11064 9222 11116 9274
rect 5448 9120 5500 9172
rect 6644 9120 6696 9172
rect 9588 9120 9640 9172
rect 9680 9120 9732 9172
rect 11336 9120 11388 9172
rect 9956 9052 10008 9104
rect 1768 8984 1820 9036
rect 8484 8984 8536 9036
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 5632 8916 5684 8968
rect 2780 8848 2832 8900
rect 5816 8959 5868 8968
rect 5816 8925 5825 8959
rect 5825 8925 5859 8959
rect 5859 8925 5868 8959
rect 5816 8916 5868 8925
rect 6000 8848 6052 8900
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 6552 8916 6604 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 6736 8848 6788 8900
rect 9680 8848 9732 8900
rect 9864 8848 9916 8900
rect 11612 8780 11664 8832
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 8894 8678 8946 8730
rect 8958 8678 9010 8730
rect 9022 8678 9074 8730
rect 9086 8678 9138 8730
rect 2136 8576 2188 8628
rect 9680 8576 9732 8628
rect 8300 8508 8352 8560
rect 9588 8483 9640 8492
rect 8116 8304 8168 8356
rect 9312 8372 9364 8424
rect 9588 8449 9597 8483
rect 9597 8449 9631 8483
rect 9631 8449 9640 8483
rect 9588 8440 9640 8449
rect 9680 8483 9732 8492
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 10692 8372 10744 8424
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 9864 8304 9916 8356
rect 2960 8134 3012 8186
rect 3024 8134 3076 8186
rect 3088 8134 3140 8186
rect 3152 8134 3204 8186
rect 6916 8134 6968 8186
rect 6980 8134 7032 8186
rect 7044 8134 7096 8186
rect 7108 8134 7160 8186
rect 10872 8134 10924 8186
rect 10936 8134 10988 8186
rect 11000 8134 11052 8186
rect 11064 8134 11116 8186
rect 3332 8032 3384 8084
rect 2596 7964 2648 8016
rect 2872 7964 2924 8016
rect 6736 7964 6788 8016
rect 7840 7964 7892 8016
rect 3240 7896 3292 7948
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 3516 7828 3568 7880
rect 7840 7828 7892 7880
rect 12256 7871 12308 7880
rect 12256 7837 12265 7871
rect 12265 7837 12299 7871
rect 12299 7837 12308 7871
rect 12256 7828 12308 7837
rect 1492 7735 1544 7744
rect 1492 7701 1501 7735
rect 1501 7701 1535 7735
rect 1535 7701 1544 7735
rect 1492 7692 1544 7701
rect 2504 7735 2556 7744
rect 2504 7701 2513 7735
rect 2513 7701 2547 7735
rect 2547 7701 2556 7735
rect 2504 7692 2556 7701
rect 2688 7760 2740 7812
rect 9680 7760 9732 7812
rect 3516 7692 3568 7744
rect 3976 7692 4028 7744
rect 6460 7692 6512 7744
rect 8024 7692 8076 7744
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 8894 7590 8946 7642
rect 8958 7590 9010 7642
rect 9022 7590 9074 7642
rect 9086 7590 9138 7642
rect 6460 7488 6512 7540
rect 7656 7488 7708 7540
rect 2136 7352 2188 7404
rect 7288 7420 7340 7472
rect 2504 7352 2556 7404
rect 3240 7352 3292 7404
rect 3424 7352 3476 7404
rect 11428 7352 11480 7404
rect 2688 7284 2740 7336
rect 2780 7284 2832 7336
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8024 7284 8076 7336
rect 8300 7284 8352 7336
rect 7472 7216 7524 7268
rect 9588 7216 9640 7268
rect 8024 7148 8076 7200
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 2960 7046 3012 7098
rect 3024 7046 3076 7098
rect 3088 7046 3140 7098
rect 3152 7046 3204 7098
rect 6916 7046 6968 7098
rect 6980 7046 7032 7098
rect 7044 7046 7096 7098
rect 7108 7046 7160 7098
rect 10872 7046 10924 7098
rect 10936 7046 10988 7098
rect 11000 7046 11052 7098
rect 11064 7046 11116 7098
rect 2136 6944 2188 6996
rect 6736 6944 6788 6996
rect 7472 6944 7524 6996
rect 7748 6944 7800 6996
rect 3424 6876 3476 6928
rect 6368 6876 6420 6928
rect 2872 6808 2924 6860
rect 5540 6808 5592 6860
rect 6276 6808 6328 6860
rect 2228 6783 2280 6792
rect 2228 6749 2237 6783
rect 2237 6749 2271 6783
rect 2271 6749 2280 6783
rect 2228 6740 2280 6749
rect 2688 6740 2740 6792
rect 4252 6740 4304 6792
rect 4528 6740 4580 6792
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 7012 6876 7064 6928
rect 7196 6876 7248 6928
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 7472 6808 7524 6860
rect 8392 6808 8444 6860
rect 7656 6740 7708 6792
rect 6092 6672 6144 6724
rect 1584 6604 1636 6656
rect 3608 6604 3660 6656
rect 3976 6604 4028 6656
rect 4160 6604 4212 6656
rect 7104 6672 7156 6724
rect 9220 6808 9272 6860
rect 8576 6740 8628 6792
rect 12164 6808 12216 6860
rect 8852 6672 8904 6724
rect 9496 6604 9548 6656
rect 10140 6672 10192 6724
rect 10784 6672 10836 6724
rect 12072 6715 12124 6724
rect 12072 6681 12081 6715
rect 12081 6681 12115 6715
rect 12115 6681 12124 6715
rect 12072 6672 12124 6681
rect 10232 6604 10284 6656
rect 12164 6647 12216 6656
rect 12164 6613 12173 6647
rect 12173 6613 12207 6647
rect 12207 6613 12216 6647
rect 12164 6604 12216 6613
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 8894 6502 8946 6554
rect 8958 6502 9010 6554
rect 9022 6502 9074 6554
rect 9086 6502 9138 6554
rect 3332 6400 3384 6452
rect 5356 6400 5408 6452
rect 6368 6400 6420 6452
rect 8208 6400 8260 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2688 6264 2740 6316
rect 2872 6307 2924 6316
rect 2872 6273 2881 6307
rect 2881 6273 2915 6307
rect 2915 6273 2924 6307
rect 2872 6264 2924 6273
rect 4068 6264 4120 6316
rect 7196 6332 7248 6384
rect 9864 6400 9916 6452
rect 10232 6400 10284 6452
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 6092 6264 6144 6316
rect 6644 6264 6696 6316
rect 7012 6264 7064 6316
rect 7656 6264 7708 6316
rect 8300 6264 8352 6316
rect 9220 6307 9272 6316
rect 9220 6273 9229 6307
rect 9229 6273 9263 6307
rect 9263 6273 9272 6307
rect 9220 6264 9272 6273
rect 9588 6264 9640 6316
rect 9772 6264 9824 6316
rect 10416 6307 10468 6316
rect 10416 6273 10425 6307
rect 10425 6273 10459 6307
rect 10459 6273 10468 6307
rect 10416 6264 10468 6273
rect 9404 6196 9456 6248
rect 10048 6196 10100 6248
rect 11244 6196 11296 6248
rect 11520 6196 11572 6248
rect 2780 6128 2832 6180
rect 2688 6060 2740 6112
rect 8760 6128 8812 6180
rect 9036 6128 9088 6180
rect 9772 6128 9824 6180
rect 10784 6128 10836 6180
rect 3608 6060 3660 6112
rect 4804 6060 4856 6112
rect 5356 6060 5408 6112
rect 6736 6060 6788 6112
rect 2960 5958 3012 6010
rect 3024 5958 3076 6010
rect 3088 5958 3140 6010
rect 3152 5958 3204 6010
rect 6916 5958 6968 6010
rect 6980 5958 7032 6010
rect 7044 5958 7096 6010
rect 7108 5958 7160 6010
rect 10872 5958 10924 6010
rect 10936 5958 10988 6010
rect 11000 5958 11052 6010
rect 11064 5958 11116 6010
rect 4528 5763 4580 5772
rect 4528 5729 4537 5763
rect 4537 5729 4571 5763
rect 4571 5729 4580 5763
rect 4528 5720 4580 5729
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 7288 5856 7340 5908
rect 7656 5856 7708 5908
rect 10416 5856 10468 5908
rect 11704 5856 11756 5908
rect 5724 5788 5776 5840
rect 6644 5720 6696 5772
rect 6828 5720 6880 5772
rect 5908 5652 5960 5704
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 9128 5720 9180 5772
rect 9588 5720 9640 5772
rect 7656 5584 7708 5636
rect 10140 5652 10192 5704
rect 10232 5584 10284 5636
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 5540 5516 5592 5568
rect 8300 5516 8352 5568
rect 11980 5720 12032 5772
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10876 5695 10928 5704
rect 10600 5652 10652 5661
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11244 5652 11296 5704
rect 10784 5584 10836 5636
rect 11980 5627 12032 5636
rect 11980 5593 11989 5627
rect 11989 5593 12023 5627
rect 12023 5593 12032 5627
rect 11980 5584 12032 5593
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 8894 5414 8946 5466
rect 8958 5414 9010 5466
rect 9022 5414 9074 5466
rect 9086 5414 9138 5466
rect 5816 5312 5868 5364
rect 5908 5312 5960 5364
rect 7932 5312 7984 5364
rect 7472 5244 7524 5296
rect 10600 5244 10652 5296
rect 10876 5244 10928 5296
rect 11888 5287 11940 5296
rect 11888 5253 11897 5287
rect 11897 5253 11931 5287
rect 11931 5253 11940 5287
rect 11888 5244 11940 5253
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 4160 5176 4212 5228
rect 5816 5176 5868 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 7840 5176 7892 5228
rect 11244 5176 11296 5228
rect 5908 5108 5960 5160
rect 9220 5108 9272 5160
rect 10324 5040 10376 5092
rect 11244 5040 11296 5092
rect 11980 5040 12032 5092
rect 4528 4972 4580 5024
rect 2960 4870 3012 4922
rect 3024 4870 3076 4922
rect 3088 4870 3140 4922
rect 3152 4870 3204 4922
rect 6916 4870 6968 4922
rect 6980 4870 7032 4922
rect 7044 4870 7096 4922
rect 7108 4870 7160 4922
rect 10872 4870 10924 4922
rect 10936 4870 10988 4922
rect 11000 4870 11052 4922
rect 11064 4870 11116 4922
rect 2228 4768 2280 4820
rect 4620 4768 4672 4820
rect 5540 4768 5592 4820
rect 5908 4768 5960 4820
rect 8392 4768 8444 4820
rect 6000 4700 6052 4752
rect 3608 4632 3660 4684
rect 8484 4632 8536 4684
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 3884 4564 3936 4616
rect 3976 4428 4028 4480
rect 4252 4564 4304 4616
rect 6644 4564 6696 4616
rect 8208 4564 8260 4616
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 7288 4496 7340 4548
rect 11520 4539 11572 4548
rect 11520 4505 11529 4539
rect 11529 4505 11563 4539
rect 11563 4505 11572 4539
rect 11520 4496 11572 4505
rect 5264 4428 5316 4480
rect 8392 4428 8444 4480
rect 11888 4428 11940 4480
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 8894 4326 8946 4378
rect 8958 4326 9010 4378
rect 9022 4326 9074 4378
rect 9086 4326 9138 4378
rect 2780 4224 2832 4276
rect 4712 4224 4764 4276
rect 8392 4224 8444 4276
rect 8668 4224 8720 4276
rect 8300 4156 8352 4208
rect 5356 4088 5408 4140
rect 7748 4088 7800 4140
rect 8392 4020 8444 4072
rect 10324 4088 10376 4140
rect 10508 4088 10560 4140
rect 9496 4020 9548 4072
rect 11888 4199 11940 4208
rect 11888 4165 11897 4199
rect 11897 4165 11931 4199
rect 11931 4165 11940 4199
rect 11888 4156 11940 4165
rect 7472 3952 7524 4004
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 9404 3952 9456 4004
rect 9956 3995 10008 4004
rect 9956 3961 9965 3995
rect 9965 3961 9999 3995
rect 9999 3961 10008 3995
rect 9956 3952 10008 3961
rect 11796 4020 11848 4072
rect 10692 3884 10744 3936
rect 2960 3782 3012 3834
rect 3024 3782 3076 3834
rect 3088 3782 3140 3834
rect 3152 3782 3204 3834
rect 6916 3782 6968 3834
rect 6980 3782 7032 3834
rect 7044 3782 7096 3834
rect 7108 3782 7160 3834
rect 10872 3782 10924 3834
rect 10936 3782 10988 3834
rect 11000 3782 11052 3834
rect 11064 3782 11116 3834
rect 5632 3680 5684 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 10416 3680 10468 3732
rect 6460 3612 6512 3664
rect 9312 3544 9364 3596
rect 9496 3544 9548 3596
rect 11980 3587 12032 3596
rect 11980 3553 11989 3587
rect 11989 3553 12023 3587
rect 12023 3553 12032 3587
rect 11980 3544 12032 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 5724 3408 5776 3460
rect 10048 3476 10100 3528
rect 12900 3476 12952 3528
rect 10508 3408 10560 3460
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 8894 3238 8946 3290
rect 8958 3238 9010 3290
rect 9022 3238 9074 3290
rect 9086 3238 9138 3290
rect 7288 3136 7340 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 12164 3179 12216 3188
rect 9680 3136 9732 3145
rect 12164 3145 12173 3179
rect 12173 3145 12207 3179
rect 12207 3145 12216 3179
rect 12164 3136 12216 3145
rect 6276 3068 6328 3120
rect 20 3000 72 3052
rect 10600 3068 10652 3120
rect 8852 3000 8904 3052
rect 11336 3068 11388 3120
rect 9220 2864 9272 2916
rect 3700 2796 3752 2848
rect 2960 2694 3012 2746
rect 3024 2694 3076 2746
rect 3088 2694 3140 2746
rect 3152 2694 3204 2746
rect 6916 2694 6968 2746
rect 6980 2694 7032 2746
rect 7044 2694 7096 2746
rect 7108 2694 7160 2746
rect 10872 2694 10924 2746
rect 10936 2694 10988 2746
rect 11000 2694 11052 2746
rect 11064 2694 11116 2746
rect 6552 2524 6604 2576
rect 7380 2524 7432 2576
rect 8576 2524 8628 2576
rect 3884 2388 3936 2440
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 1308 2320 1360 2372
rect 2596 2320 2648 2372
rect 5264 2363 5316 2372
rect 5264 2329 5273 2363
rect 5273 2329 5307 2363
rect 5307 2329 5316 2363
rect 5264 2320 5316 2329
rect 6460 2388 6512 2440
rect 9680 2456 9732 2508
rect 11428 2592 11480 2644
rect 11612 2592 11664 2644
rect 11520 2524 11572 2576
rect 8024 2431 8076 2440
rect 8024 2397 8033 2431
rect 8033 2397 8067 2431
rect 8067 2397 8076 2431
rect 8024 2388 8076 2397
rect 9220 2388 9272 2440
rect 10416 2388 10468 2440
rect 11520 2388 11572 2440
rect 7472 2252 7524 2304
rect 7748 2320 7800 2372
rect 8116 2252 8168 2304
rect 10140 2295 10192 2304
rect 10140 2261 10149 2295
rect 10149 2261 10183 2295
rect 10183 2261 10192 2295
rect 10140 2252 10192 2261
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 8894 2150 8946 2202
rect 8958 2150 9010 2202
rect 9022 2150 9074 2202
rect 9086 2150 9138 2202
rect 9588 2048 9640 2100
rect 10140 2048 10192 2100
<< metal2 >>
rect 570 15506 626 16306
rect 1858 15506 1914 16306
rect 3146 15506 3202 16306
rect 3252 15558 3464 15586
rect 584 12918 612 15506
rect 1766 13424 1822 13433
rect 1872 13394 1900 15506
rect 3160 15450 3188 15506
rect 3252 15450 3280 15558
rect 3160 15422 3280 15450
rect 2778 15328 2834 15337
rect 2778 15263 2834 15272
rect 1766 13359 1768 13368
rect 1820 13359 1822 13368
rect 1860 13388 1912 13394
rect 1768 13330 1820 13336
rect 1860 13330 1912 13336
rect 2792 13326 2820 15263
rect 2934 13628 3230 13648
rect 2990 13626 3014 13628
rect 3070 13626 3094 13628
rect 3150 13626 3174 13628
rect 3012 13574 3014 13626
rect 3076 13574 3088 13626
rect 3150 13574 3152 13626
rect 2990 13572 3014 13574
rect 3070 13572 3094 13574
rect 3150 13572 3174 13574
rect 2934 13552 3230 13572
rect 3436 13462 3464 15558
rect 4434 15506 4490 16306
rect 5722 15506 5778 16306
rect 7010 15506 7066 16306
rect 7116 15558 7328 15586
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 4448 13326 4476 15506
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 572 12912 624 12918
rect 572 12854 624 12860
rect 1504 12434 1532 13194
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 2700 12986 2728 13126
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 3976 12912 4028 12918
rect 4028 12860 4384 12866
rect 3976 12854 4384 12860
rect 3988 12850 4384 12854
rect 3424 12844 3476 12850
rect 3424 12786 3476 12792
rect 3988 12844 4396 12850
rect 3988 12838 4344 12844
rect 2934 12540 3230 12560
rect 2990 12538 3014 12540
rect 3070 12538 3094 12540
rect 3150 12538 3174 12540
rect 3012 12486 3014 12538
rect 3076 12486 3088 12538
rect 3150 12486 3152 12538
rect 2990 12484 3014 12486
rect 3070 12484 3094 12486
rect 3150 12484 3174 12486
rect 2934 12464 3230 12484
rect 3436 12434 3464 12786
rect 3884 12436 3936 12442
rect 1504 12406 1624 12434
rect 3436 12406 3556 12434
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 11529 1440 11630
rect 1398 11520 1454 11529
rect 1398 11455 1454 11464
rect 1492 7744 1544 7750
rect 1490 7712 1492 7721
rect 1544 7712 1546 7721
rect 1490 7647 1546 7656
rect 1596 6662 1624 12406
rect 1768 12164 1820 12170
rect 1768 12106 1820 12112
rect 1780 9042 1808 12106
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1872 9625 1900 9930
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9722 1992 9862
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1858 9616 1914 9625
rect 1858 9551 1914 9560
rect 1768 9036 1820 9042
rect 1768 8978 1820 8984
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8634 2176 8910
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 7002 2176 7346
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2228 6792 2280 6798
rect 2424 6769 2452 12038
rect 2934 11452 3230 11472
rect 2990 11450 3014 11452
rect 3070 11450 3094 11452
rect 3150 11450 3174 11452
rect 3012 11398 3014 11450
rect 3076 11398 3088 11450
rect 3150 11398 3152 11450
rect 2990 11396 3014 11398
rect 3070 11396 3094 11398
rect 3150 11396 3174 11398
rect 2934 11376 3230 11396
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 2934 10364 3230 10384
rect 2990 10362 3014 10364
rect 3070 10362 3094 10364
rect 3150 10362 3174 10364
rect 3012 10310 3014 10362
rect 3076 10310 3088 10362
rect 3150 10310 3152 10362
rect 2990 10308 3014 10310
rect 3070 10308 3094 10310
rect 3150 10308 3174 10310
rect 2934 10288 3230 10308
rect 3332 10192 3384 10198
rect 3332 10134 3384 10140
rect 2934 9276 3230 9296
rect 2990 9274 3014 9276
rect 3070 9274 3094 9276
rect 3150 9274 3174 9276
rect 3012 9222 3014 9274
rect 3076 9222 3088 9274
rect 3150 9222 3152 9274
rect 2990 9220 3014 9222
rect 3070 9220 3094 9222
rect 3150 9220 3174 9222
rect 2934 9200 3230 9220
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2608 7834 2636 7958
rect 2608 7818 2728 7834
rect 2608 7812 2740 7818
rect 2608 7806 2688 7812
rect 2688 7754 2740 7760
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7410 2544 7686
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2792 7342 2820 8842
rect 2934 8188 3230 8208
rect 2990 8186 3014 8188
rect 3070 8186 3094 8188
rect 3150 8186 3174 8188
rect 3012 8134 3014 8186
rect 3076 8134 3088 8186
rect 3150 8134 3152 8186
rect 2990 8132 3014 8134
rect 3070 8132 3094 8134
rect 3150 8132 3174 8134
rect 2934 8112 3230 8132
rect 3344 8090 3372 10134
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2700 6798 2728 7278
rect 2884 7188 2912 7958
rect 3240 7948 3292 7954
rect 3436 7936 3464 11086
rect 3240 7890 3292 7896
rect 3344 7908 3464 7936
rect 3252 7410 3280 7890
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 2792 7160 2912 7188
rect 2688 6792 2740 6798
rect 2228 6734 2280 6740
rect 2410 6760 2466 6769
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5817 1440 6258
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 2240 4826 2268 6734
rect 2688 6734 2740 6740
rect 2410 6695 2466 6704
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 6118 2728 6258
rect 2792 6186 2820 7160
rect 2934 7100 3230 7120
rect 2990 7098 3014 7100
rect 3070 7098 3094 7100
rect 3150 7098 3174 7100
rect 3012 7046 3014 7098
rect 3076 7046 3088 7098
rect 3150 7046 3152 7098
rect 2990 7044 3014 7046
rect 3070 7044 3094 7046
rect 3150 7044 3174 7046
rect 2934 7024 3230 7044
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 2884 6322 2912 6802
rect 3344 6458 3372 7908
rect 3528 7886 3556 12406
rect 3988 12434 4016 12838
rect 4344 12786 4396 12792
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3988 12406 4108 12434
rect 3884 12378 3936 12384
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3436 6934 3464 7346
rect 3424 6928 3476 6934
rect 3424 6870 3476 6876
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2792 4282 2820 6122
rect 2934 6012 3230 6032
rect 2990 6010 3014 6012
rect 3070 6010 3094 6012
rect 3150 6010 3174 6012
rect 3012 5958 3014 6010
rect 3076 5958 3088 6010
rect 3150 5958 3152 6010
rect 2990 5956 3014 5958
rect 3070 5956 3094 5958
rect 3150 5956 3174 5958
rect 2934 5936 3230 5956
rect 3436 5234 3464 6870
rect 3528 5234 3556 7686
rect 3620 6662 3648 11494
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 2934 4924 3230 4944
rect 2990 4922 3014 4924
rect 3070 4922 3094 4924
rect 3150 4922 3174 4924
rect 3012 4870 3014 4922
rect 3076 4870 3088 4922
rect 3150 4870 3152 4922
rect 2990 4868 3014 4870
rect 3070 4868 3094 4870
rect 3150 4868 3174 4870
rect 2934 4848 3230 4868
rect 3620 4690 3648 6054
rect 3608 4684 3660 4690
rect 3608 4626 3660 4632
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 1860 3936 1912 3942
rect 1858 3904 1860 3913
rect 1912 3904 1914 3913
rect 1858 3839 1914 3848
rect 2934 3836 3230 3856
rect 2990 3834 3014 3836
rect 3070 3834 3094 3836
rect 3150 3834 3174 3836
rect 3012 3782 3014 3834
rect 3076 3782 3088 3834
rect 3150 3782 3152 3834
rect 2990 3780 3014 3782
rect 3070 3780 3094 3782
rect 3150 3780 3174 3782
rect 2934 3760 3230 3780
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 20 3052 72 3058
rect 20 2994 72 3000
rect 32 800 60 2994
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 800 1348 2314
rect 1412 2009 1440 3470
rect 3712 2854 3740 12310
rect 3792 12232 3844 12238
rect 3790 12200 3792 12209
rect 3844 12200 3846 12209
rect 3790 12135 3846 12144
rect 3896 11558 3924 12378
rect 4080 12238 4108 12406
rect 4172 12306 4200 12582
rect 4160 12300 4212 12306
rect 4160 12242 4212 12248
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3804 10266 3832 11018
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3804 4622 3832 10202
rect 3896 4622 3924 11222
rect 3988 7750 4016 11494
rect 4080 11150 4108 12174
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 3988 4486 4016 6598
rect 4080 6322 4108 9862
rect 4264 6798 4292 12650
rect 4344 12232 4396 12238
rect 4342 12200 4344 12209
rect 4396 12200 4398 12209
rect 4448 12170 4476 12718
rect 4342 12135 4398 12144
rect 4436 12164 4488 12170
rect 4436 12106 4488 12112
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4356 10062 4384 10202
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4172 5234 4200 6598
rect 4356 6474 4384 9998
rect 4264 6446 4384 6474
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4264 4622 4292 6446
rect 4448 6361 4476 12106
rect 4540 10062 4568 13126
rect 4912 13084 5208 13104
rect 4968 13082 4992 13084
rect 5048 13082 5072 13084
rect 5128 13082 5152 13084
rect 4990 13030 4992 13082
rect 5054 13030 5066 13082
rect 5128 13030 5130 13082
rect 4968 13028 4992 13030
rect 5048 13028 5072 13030
rect 5128 13028 5152 13030
rect 4912 13008 5208 13028
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4434 6352 4490 6361
rect 4434 6287 4490 6296
rect 4434 6216 4490 6225
rect 4434 6151 4490 6160
rect 4448 5710 4476 6151
rect 4540 5778 4568 6734
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4540 5030 4568 5714
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4632 4826 4660 12854
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4724 12434 4752 12786
rect 4724 12406 4844 12434
rect 4710 11656 4766 11665
rect 4710 11591 4766 11600
rect 4724 11354 4752 11591
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4724 10742 4752 11154
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 4724 4282 4752 10678
rect 4816 6118 4844 12406
rect 4912 11996 5208 12016
rect 4968 11994 4992 11996
rect 5048 11994 5072 11996
rect 5128 11994 5152 11996
rect 4990 11942 4992 11994
rect 5054 11942 5066 11994
rect 5128 11942 5130 11994
rect 4968 11940 4992 11942
rect 5048 11940 5072 11942
rect 5128 11940 5152 11942
rect 4912 11920 5208 11940
rect 5276 11218 5304 13126
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 4912 10908 5208 10928
rect 4968 10906 4992 10908
rect 5048 10906 5072 10908
rect 5128 10906 5152 10908
rect 4990 10854 4992 10906
rect 5054 10854 5066 10906
rect 5128 10854 5130 10906
rect 4968 10852 4992 10854
rect 5048 10852 5072 10854
rect 5128 10852 5152 10854
rect 4912 10832 5208 10852
rect 4912 9820 5208 9840
rect 4968 9818 4992 9820
rect 5048 9818 5072 9820
rect 5128 9818 5152 9820
rect 4990 9766 4992 9818
rect 5054 9766 5066 9818
rect 5128 9766 5130 9818
rect 4968 9764 4992 9766
rect 5048 9764 5072 9766
rect 5128 9764 5152 9766
rect 4912 9744 5208 9764
rect 4912 8732 5208 8752
rect 4968 8730 4992 8732
rect 5048 8730 5072 8732
rect 5128 8730 5152 8732
rect 4990 8678 4992 8730
rect 5054 8678 5066 8730
rect 5128 8678 5130 8730
rect 4968 8676 4992 8678
rect 5048 8676 5072 8678
rect 5128 8676 5152 8678
rect 4912 8656 5208 8676
rect 4912 7644 5208 7664
rect 4968 7642 4992 7644
rect 5048 7642 5072 7644
rect 5128 7642 5152 7644
rect 4990 7590 4992 7642
rect 5054 7590 5066 7642
rect 5128 7590 5130 7642
rect 4968 7588 4992 7590
rect 5048 7588 5072 7590
rect 5128 7588 5152 7590
rect 4912 7568 5208 7588
rect 4912 6556 5208 6576
rect 4968 6554 4992 6556
rect 5048 6554 5072 6556
rect 5128 6554 5152 6556
rect 4990 6502 4992 6554
rect 5054 6502 5066 6554
rect 5128 6502 5130 6554
rect 4968 6500 4992 6502
rect 5048 6500 5072 6502
rect 5128 6500 5152 6502
rect 4912 6480 5208 6500
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4912 5468 5208 5488
rect 4968 5466 4992 5468
rect 5048 5466 5072 5468
rect 5128 5466 5152 5468
rect 4990 5414 4992 5466
rect 5054 5414 5066 5466
rect 5128 5414 5130 5466
rect 4968 5412 4992 5414
rect 5048 5412 5072 5414
rect 5128 5412 5152 5414
rect 4912 5392 5208 5412
rect 5276 4486 5304 10950
rect 5368 6458 5396 13466
rect 5736 13462 5764 15506
rect 7024 15450 7052 15506
rect 7116 15450 7144 15558
rect 7024 15422 7144 15450
rect 6890 13628 7186 13648
rect 6946 13626 6970 13628
rect 7026 13626 7050 13628
rect 7106 13626 7130 13628
rect 6968 13574 6970 13626
rect 7032 13574 7044 13626
rect 7106 13574 7108 13626
rect 6946 13572 6970 13574
rect 7026 13572 7050 13574
rect 7106 13572 7130 13574
rect 6890 13552 7186 13572
rect 7300 13462 7328 15558
rect 8298 15506 8354 16306
rect 9232 15558 9536 15586
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5460 9178 5488 13194
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5552 10810 5580 12854
rect 6564 12434 6592 13126
rect 7288 12708 7340 12714
rect 7288 12650 7340 12656
rect 6890 12540 7186 12560
rect 6946 12538 6970 12540
rect 7026 12538 7050 12540
rect 7106 12538 7130 12540
rect 6968 12486 6970 12538
rect 7032 12486 7044 12538
rect 7106 12486 7108 12538
rect 6946 12484 6970 12486
rect 7026 12484 7050 12486
rect 7106 12484 7130 12486
rect 6890 12464 7186 12484
rect 6564 12406 6684 12434
rect 6000 12232 6052 12238
rect 6000 12174 6052 12180
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5552 8922 5580 9862
rect 5460 8894 5580 8922
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 6118 5396 6394
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5460 5930 5488 8894
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 6866 5580 8774
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5368 5902 5488 5930
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 4912 4380 5208 4400
rect 4968 4378 4992 4380
rect 5048 4378 5072 4380
rect 5128 4378 5152 4380
rect 4990 4326 4992 4378
rect 5054 4326 5066 4378
rect 5128 4326 5130 4378
rect 4968 4324 4992 4326
rect 5048 4324 5072 4326
rect 5128 4324 5152 4326
rect 4912 4304 5208 4324
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 5368 4146 5396 5902
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 4912 3292 5208 3312
rect 4968 3290 4992 3292
rect 5048 3290 5072 3292
rect 5128 3290 5152 3292
rect 4990 3238 4992 3290
rect 5054 3238 5066 3290
rect 5128 3238 5130 3290
rect 4968 3236 4992 3238
rect 5048 3236 5072 3238
rect 5128 3236 5152 3238
rect 4912 3216 5208 3236
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 2934 2748 3230 2768
rect 2990 2746 3014 2748
rect 3070 2746 3094 2748
rect 3150 2746 3174 2748
rect 3012 2694 3014 2746
rect 3076 2694 3088 2746
rect 3150 2694 3152 2746
rect 2990 2692 3014 2694
rect 3070 2692 3094 2694
rect 3150 2692 3174 2694
rect 2934 2672 3230 2692
rect 5460 2446 5488 5510
rect 5552 4826 5580 5510
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5644 3738 5672 8910
rect 5736 5846 5764 11630
rect 5828 8974 5856 12038
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5736 3466 5764 5782
rect 5828 5370 5856 8910
rect 6012 8906 6040 12174
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 10810 6408 11698
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 11150 6500 11562
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5370 5948 5646
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5814 5264 5870 5273
rect 5814 5199 5816 5208
rect 5868 5199 5870 5208
rect 5816 5170 5868 5176
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 4826 5948 5102
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6012 4758 6040 8842
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6104 6322 6132 6666
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6196 5710 6224 10474
rect 6288 9722 6316 10474
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6380 6934 6408 9658
rect 6656 9586 6684 12406
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6932 11665 6960 11698
rect 6918 11656 6974 11665
rect 6918 11591 6974 11600
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6656 9178 6684 9522
rect 6748 9382 6776 11494
rect 6890 11452 7186 11472
rect 6946 11450 6970 11452
rect 7026 11450 7050 11452
rect 7106 11450 7130 11452
rect 6968 11398 6970 11450
rect 7032 11398 7044 11450
rect 7106 11398 7108 11450
rect 6946 11396 6970 11398
rect 7026 11396 7050 11398
rect 7106 11396 7130 11398
rect 6890 11376 7186 11396
rect 7300 11234 7328 12650
rect 7300 11206 7420 11234
rect 7288 11076 7340 11082
rect 7288 11018 7340 11024
rect 6890 10364 7186 10384
rect 6946 10362 6970 10364
rect 7026 10362 7050 10364
rect 7106 10362 7130 10364
rect 6968 10310 6970 10362
rect 7032 10310 7044 10362
rect 7106 10310 7108 10362
rect 6946 10308 6970 10310
rect 7026 10308 7050 10310
rect 7106 10308 7130 10310
rect 6890 10288 7186 10308
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6472 7546 6500 7686
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 6928 6420 6934
rect 6420 6876 6500 6882
rect 6368 6870 6500 6876
rect 6276 6860 6328 6866
rect 6380 6854 6500 6870
rect 6276 6802 6328 6808
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 6288 3126 6316 6802
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6380 6458 6408 6734
rect 6368 6452 6420 6458
rect 6368 6394 6420 6400
rect 6472 3670 6500 6854
rect 6564 5234 6592 8910
rect 6748 8906 6776 9318
rect 6890 9276 7186 9296
rect 6946 9274 6970 9276
rect 7026 9274 7050 9276
rect 7106 9274 7130 9276
rect 6968 9222 6970 9274
rect 7032 9222 7044 9274
rect 7106 9222 7108 9274
rect 6946 9220 6970 9222
rect 7026 9220 7050 9222
rect 7106 9220 7130 9222
rect 6890 9200 7186 9220
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6890 8188 7186 8208
rect 6946 8186 6970 8188
rect 7026 8186 7050 8188
rect 7106 8186 7130 8188
rect 6968 8134 6970 8186
rect 7032 8134 7044 8186
rect 7106 8134 7108 8186
rect 6946 8132 6970 8134
rect 7026 8132 7050 8134
rect 7106 8132 7130 8134
rect 6890 8112 7186 8132
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6748 7002 6776 7958
rect 7300 7478 7328 11018
rect 7392 10470 7420 11206
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7484 10266 7512 13126
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 7576 11218 7604 12650
rect 8036 12434 8064 13670
rect 8312 13326 8340 15506
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12850 8340 13126
rect 8868 13084 9164 13104
rect 8924 13082 8948 13084
rect 9004 13082 9028 13084
rect 9084 13082 9108 13084
rect 8946 13030 8948 13082
rect 9010 13030 9022 13082
rect 9084 13030 9086 13082
rect 8924 13028 8948 13030
rect 9004 13028 9028 13030
rect 9084 13028 9108 13030
rect 8868 13008 9164 13028
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 7852 12406 8064 12434
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7288 7472 7340 7478
rect 7288 7414 7340 7420
rect 6890 7100 7186 7120
rect 6946 7098 6970 7100
rect 7026 7098 7050 7100
rect 7106 7098 7130 7100
rect 6968 7046 6970 7098
rect 7032 7046 7044 7098
rect 7106 7046 7108 7098
rect 6946 7044 6970 7046
rect 7026 7044 7050 7046
rect 7106 7044 7130 7046
rect 6890 7024 7186 7044
rect 6736 6996 6788 7002
rect 6736 6938 6788 6944
rect 7012 6928 7064 6934
rect 7196 6928 7248 6934
rect 7012 6870 7064 6876
rect 7102 6896 7158 6905
rect 6734 6352 6790 6361
rect 6644 6316 6696 6322
rect 7024 6322 7052 6870
rect 7196 6870 7248 6876
rect 7102 6831 7158 6840
rect 7116 6730 7144 6831
rect 7208 6798 7236 6870
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7194 6488 7250 6497
rect 7194 6423 7250 6432
rect 7208 6390 7236 6423
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 6734 6287 6790 6296
rect 7012 6316 7064 6322
rect 6644 6258 6696 6264
rect 6656 5778 6684 6258
rect 6748 6118 6776 6287
rect 7012 6258 7064 6264
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6890 6012 7186 6032
rect 6946 6010 6970 6012
rect 7026 6010 7050 6012
rect 7106 6010 7130 6012
rect 6968 5958 6970 6010
rect 7032 5958 7044 6010
rect 7106 5958 7108 6010
rect 6946 5956 6970 5958
rect 7026 5956 7050 5958
rect 7106 5956 7130 5958
rect 6890 5936 7186 5956
rect 7300 5914 7328 7414
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6826 5808 6882 5817
rect 6644 5772 6696 5778
rect 6826 5743 6828 5752
rect 6644 5714 6696 5720
rect 6880 5743 6882 5752
rect 6828 5714 6880 5720
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6564 2582 6592 5170
rect 6656 4622 6684 5714
rect 6890 4924 7186 4944
rect 6946 4922 6970 4924
rect 7026 4922 7050 4924
rect 7106 4922 7130 4924
rect 6968 4870 6970 4922
rect 7032 4870 7044 4922
rect 7106 4870 7108 4922
rect 6946 4868 6970 4870
rect 7026 4868 7050 4870
rect 7106 4868 7130 4870
rect 6890 4848 7186 4868
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 6890 3836 7186 3856
rect 6946 3834 6970 3836
rect 7026 3834 7050 3836
rect 7106 3834 7130 3836
rect 6968 3782 6970 3834
rect 7032 3782 7044 3834
rect 7106 3782 7108 3834
rect 6946 3780 6970 3782
rect 7026 3780 7050 3782
rect 7106 3780 7130 3782
rect 6890 3760 7186 3780
rect 7300 3194 7328 4490
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 6890 2748 7186 2768
rect 6946 2746 6970 2748
rect 7026 2746 7050 2748
rect 7106 2746 7130 2748
rect 6968 2694 6970 2746
rect 7032 2694 7044 2746
rect 7106 2694 7108 2746
rect 6946 2692 6970 2694
rect 7026 2692 7050 2694
rect 7106 2692 7130 2694
rect 6890 2672 7186 2692
rect 7392 2582 7420 9318
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7484 7002 7512 7210
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7484 5302 7512 6802
rect 7576 5760 7604 10406
rect 7668 7546 7696 12038
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7668 6798 7696 7482
rect 7760 7177 7788 10678
rect 7852 8022 7880 12406
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8404 11762 8432 12242
rect 9232 12238 9260 15558
rect 9508 15450 9536 15558
rect 9586 15506 9642 16306
rect 10874 15506 10930 16306
rect 12162 15506 12218 16306
rect 13450 15506 13506 16306
rect 9600 15450 9628 15506
rect 9508 15422 9628 15450
rect 10598 15328 10654 15337
rect 10598 15263 10654 15272
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 13326 9812 13670
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9600 13138 9628 13194
rect 9600 13110 10180 13138
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 8868 11996 9164 12016
rect 8924 11994 8948 11996
rect 9004 11994 9028 11996
rect 9084 11994 9108 11996
rect 8946 11942 8948 11994
rect 9010 11942 9022 11994
rect 9084 11942 9086 11994
rect 8924 11940 8948 11942
rect 9004 11940 9028 11942
rect 9084 11940 9108 11942
rect 8868 11920 9164 11940
rect 9324 11898 9352 12786
rect 9784 12434 9812 12786
rect 9692 12406 9812 12434
rect 9496 12300 9548 12306
rect 9496 12242 9548 12248
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7840 8016 7892 8022
rect 7840 7958 7892 7964
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7746 7168 7802 7177
rect 7746 7103 7802 7112
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 5914 7696 6258
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7576 5732 7696 5760
rect 7562 5672 7618 5681
rect 7668 5642 7696 5732
rect 7562 5607 7618 5616
rect 7656 5636 7708 5642
rect 7472 5296 7524 5302
rect 7472 5238 7524 5244
rect 7484 4010 7512 5238
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 7576 2774 7604 5607
rect 7656 5578 7708 5584
rect 7760 4146 7788 6938
rect 7852 5234 7880 7822
rect 8036 7750 8064 11630
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8116 8356 8168 8362
rect 8116 8298 8168 8304
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7342 8064 7686
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 7944 5370 7972 7278
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7484 2746 7604 2774
rect 6552 2576 6604 2582
rect 6552 2518 6604 2524
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 6460 2440 6512 2446
rect 6460 2382 6512 2388
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 1398 2000 1454 2009
rect 1398 1935 1454 1944
rect 2608 800 2636 2314
rect 3896 800 3924 2382
rect 5264 2372 5316 2378
rect 5264 2314 5316 2320
rect 4912 2204 5208 2224
rect 4968 2202 4992 2204
rect 5048 2202 5072 2204
rect 5128 2202 5152 2204
rect 4990 2150 4992 2202
rect 5054 2150 5066 2202
rect 5128 2150 5130 2202
rect 4968 2148 4992 2150
rect 5048 2148 5072 2150
rect 5128 2148 5152 2150
rect 4912 2128 5208 2148
rect 5276 1170 5304 2314
rect 5184 1142 5304 1170
rect 5184 800 5212 1142
rect 6472 800 6500 2382
rect 7484 2310 7512 2746
rect 8036 2446 8064 7142
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7760 800 7788 2314
rect 8128 2310 8156 8298
rect 8220 6458 8248 11018
rect 8312 8566 8340 11698
rect 9220 11552 9272 11558
rect 9220 11494 9272 11500
rect 9232 11286 9260 11494
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 8868 10908 9164 10928
rect 8924 10906 8948 10908
rect 9004 10906 9028 10908
rect 9084 10906 9108 10908
rect 8946 10854 8948 10906
rect 9010 10854 9022 10906
rect 9084 10854 9086 10906
rect 8924 10852 8948 10854
rect 9004 10852 9028 10854
rect 9084 10852 9108 10854
rect 8868 10832 9164 10852
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8220 4622 8248 6394
rect 8312 6322 8340 7278
rect 8496 7206 8524 8978
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8312 4214 8340 5510
rect 8404 4826 8432 6802
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8496 4690 8524 7142
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8588 6497 8616 6734
rect 8574 6488 8630 6497
rect 8574 6423 8630 6432
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8404 4282 8432 4422
rect 8680 4282 8708 10542
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 8772 6186 8800 9862
rect 8868 9820 9164 9840
rect 8924 9818 8948 9820
rect 9004 9818 9028 9820
rect 9084 9818 9108 9820
rect 8946 9766 8948 9818
rect 9010 9766 9022 9818
rect 9084 9766 9086 9818
rect 8924 9764 8948 9766
rect 9004 9764 9028 9766
rect 9084 9764 9108 9766
rect 8868 9744 9164 9764
rect 9324 9586 9352 11222
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9312 9376 9364 9382
rect 9312 9318 9364 9324
rect 8868 8732 9164 8752
rect 8924 8730 8948 8732
rect 9004 8730 9028 8732
rect 9084 8730 9108 8732
rect 8946 8678 8948 8730
rect 9010 8678 9022 8730
rect 9084 8678 9086 8730
rect 8924 8676 8948 8678
rect 9004 8676 9028 8678
rect 9084 8676 9108 8678
rect 8868 8656 9164 8676
rect 9324 8430 9352 9318
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9416 8362 9444 10746
rect 9508 10198 9536 12242
rect 9692 11830 9720 12406
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9496 10192 9548 10198
rect 9496 10134 9548 10140
rect 9692 9178 9720 11766
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11354 9812 11494
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9600 8498 9628 9114
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8634 9720 8842
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9784 8514 9812 11290
rect 9876 10062 9904 12922
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9968 10266 9996 12854
rect 10048 12164 10100 12170
rect 10048 12106 10100 12112
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9876 8906 9904 9998
rect 9968 9110 9996 10202
rect 10060 9450 10088 12106
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9692 8498 9812 8514
rect 9588 8492 9640 8498
rect 9588 8434 9640 8440
rect 9680 8492 9812 8498
rect 9732 8486 9812 8492
rect 9680 8434 9732 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 8868 7644 9164 7664
rect 8924 7642 8948 7644
rect 9004 7642 9028 7644
rect 9084 7642 9108 7644
rect 8946 7590 8948 7642
rect 9010 7590 9022 7642
rect 9084 7590 9086 7642
rect 8924 7588 8948 7590
rect 9004 7588 9028 7590
rect 9084 7588 9108 7590
rect 8868 7568 9164 7588
rect 8850 6896 8906 6905
rect 8850 6831 8906 6840
rect 9220 6860 9272 6866
rect 8864 6730 8892 6831
rect 9220 6802 9272 6808
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8868 6556 9164 6576
rect 8924 6554 8948 6556
rect 9004 6554 9028 6556
rect 9084 6554 9108 6556
rect 8946 6502 8948 6554
rect 9010 6502 9022 6554
rect 9084 6502 9086 6554
rect 8924 6500 8948 6502
rect 9004 6500 9028 6502
rect 9084 6500 9108 6502
rect 8868 6480 9164 6500
rect 9232 6440 9260 6802
rect 9140 6412 9260 6440
rect 9034 6216 9090 6225
rect 8760 6180 8812 6186
rect 9034 6151 9036 6160
rect 8760 6122 8812 6128
rect 9088 6151 9090 6160
rect 9036 6122 9088 6128
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8404 4078 8432 4218
rect 8392 4072 8444 4078
rect 8680 4026 8708 4218
rect 8392 4014 8444 4020
rect 8588 3998 8708 4026
rect 8588 3942 8616 3998
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8588 2582 8616 3878
rect 8772 3040 8800 6122
rect 9140 5778 9168 6412
rect 9416 6338 9444 8298
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9324 6310 9444 6338
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 8868 5468 9164 5488
rect 8924 5466 8948 5468
rect 9004 5466 9028 5468
rect 9084 5466 9108 5468
rect 8946 5414 8948 5466
rect 9010 5414 9022 5466
rect 9084 5414 9086 5466
rect 8924 5412 8948 5414
rect 9004 5412 9028 5414
rect 9084 5412 9108 5414
rect 8868 5392 9164 5412
rect 9232 5166 9260 6258
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 8868 4380 9164 4400
rect 8924 4378 8948 4380
rect 9004 4378 9028 4380
rect 9084 4378 9108 4380
rect 8946 4326 8948 4378
rect 9010 4326 9022 4378
rect 9084 4326 9086 4378
rect 8924 4324 8948 4326
rect 9004 4324 9028 4326
rect 9084 4324 9108 4326
rect 8868 4304 9164 4324
rect 8868 3292 9164 3312
rect 8924 3290 8948 3292
rect 9004 3290 9028 3292
rect 9084 3290 9108 3292
rect 8946 3238 8948 3290
rect 9010 3238 9022 3290
rect 9084 3238 9086 3290
rect 8924 3236 8948 3238
rect 9004 3236 9028 3238
rect 9084 3236 9108 3238
rect 8868 3216 9164 3236
rect 8852 3052 8904 3058
rect 8772 3012 8852 3040
rect 8852 2994 8904 3000
rect 9232 2922 9260 5102
rect 9324 3602 9352 6310
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9416 4010 9444 6190
rect 9508 4078 9536 6598
rect 9600 6322 9628 7210
rect 9692 6633 9720 7754
rect 9876 6633 9904 8298
rect 10152 6730 10180 13110
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10244 11082 10272 11290
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10244 6662 10272 9862
rect 10336 8974 10364 12650
rect 10428 11014 10456 12650
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 11008 10468 11014
rect 10416 10950 10468 10956
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10232 6656 10284 6662
rect 9678 6624 9734 6633
rect 9678 6559 9734 6568
rect 9862 6624 9918 6633
rect 10232 6598 10284 6604
rect 9862 6559 9918 6568
rect 9954 6488 10010 6497
rect 9876 6458 9954 6474
rect 9864 6452 9954 6458
rect 9916 6446 9954 6452
rect 9954 6423 10010 6432
rect 10232 6452 10284 6458
rect 9864 6394 9916 6400
rect 10232 6394 10284 6400
rect 9954 6352 10010 6361
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9772 6316 9824 6322
rect 9824 6296 9954 6304
rect 9824 6287 10010 6296
rect 9824 6276 9996 6287
rect 9772 6258 9824 6264
rect 10048 6248 10100 6254
rect 9862 6216 9918 6225
rect 9772 6180 9824 6186
rect 10244 6236 10272 6394
rect 10100 6208 10272 6236
rect 10048 6190 10100 6196
rect 9862 6151 9918 6160
rect 9772 6122 9824 6128
rect 9678 5944 9734 5953
rect 9678 5879 9734 5888
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9600 5273 9628 5714
rect 9586 5264 9642 5273
rect 9586 5199 9642 5208
rect 9496 4072 9548 4078
rect 9496 4014 9548 4020
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9508 3602 9536 4014
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 8576 2576 8628 2582
rect 8576 2518 8628 2524
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8868 2204 9164 2224
rect 8924 2202 8948 2204
rect 9004 2202 9028 2204
rect 9084 2202 9108 2204
rect 8946 2150 8948 2202
rect 9010 2150 9022 2202
rect 9084 2150 9086 2202
rect 8924 2148 8948 2150
rect 9004 2148 9028 2150
rect 9084 2148 9108 2150
rect 8868 2128 9164 2148
rect 9232 1306 9260 2382
rect 9600 2106 9628 5199
rect 9692 3194 9720 5879
rect 9784 5409 9812 6122
rect 9770 5400 9826 5409
rect 9770 5335 9826 5344
rect 9876 3738 9904 6151
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5273 10180 5646
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10244 5545 10272 5578
rect 10230 5536 10286 5545
rect 10230 5471 10286 5480
rect 10138 5264 10194 5273
rect 10138 5199 10194 5208
rect 10336 5098 10364 8910
rect 10414 6352 10470 6361
rect 10414 6287 10416 6296
rect 10468 6287 10470 6296
rect 10416 6258 10468 6264
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 9954 4040 10010 4049
rect 9954 3975 9956 3984
rect 10008 3975 10010 3984
rect 9956 3946 10008 3952
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9968 3516 9996 3946
rect 10048 3528 10100 3534
rect 9968 3488 10048 3516
rect 10048 3470 10100 3476
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9588 2100 9640 2106
rect 9588 2042 9640 2048
rect 9048 1278 9260 1306
rect 9048 800 9076 1278
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 9692 105 9720 2450
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 2106 10180 2246
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 10336 800 10364 4082
rect 10428 3738 10456 5850
rect 10520 4146 10548 12582
rect 10612 12442 10640 15263
rect 10888 13818 10916 15506
rect 10704 13790 10916 13818
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10704 11762 10732 13790
rect 10846 13628 11142 13648
rect 10902 13626 10926 13628
rect 10982 13626 11006 13628
rect 11062 13626 11086 13628
rect 10924 13574 10926 13626
rect 10988 13574 11000 13626
rect 11062 13574 11064 13626
rect 10902 13572 10926 13574
rect 10982 13572 11006 13574
rect 11062 13572 11086 13574
rect 10846 13552 11142 13572
rect 10966 13424 11022 13433
rect 10966 13359 10968 13368
rect 11020 13359 11022 13368
rect 10968 13330 11020 13336
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12986 11836 13194
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11900 12850 11928 13262
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 10846 12540 11142 12560
rect 10902 12538 10926 12540
rect 10982 12538 11006 12540
rect 11062 12538 11086 12540
rect 10924 12486 10926 12538
rect 10988 12486 11000 12538
rect 11062 12486 11064 12538
rect 10902 12484 10926 12486
rect 10982 12484 11006 12486
rect 11062 12484 11086 12486
rect 10846 12464 11142 12484
rect 11716 12434 11744 12786
rect 11992 12646 12020 12922
rect 12084 12730 12112 13194
rect 12176 12918 12204 15506
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12084 12702 12204 12730
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11716 12406 11928 12434
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 11762 10824 12310
rect 10692 11756 10744 11762
rect 10692 11698 10744 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 10846 11452 11142 11472
rect 10902 11450 10926 11452
rect 10982 11450 11006 11452
rect 11062 11450 11086 11452
rect 10924 11398 10926 11450
rect 10988 11398 11000 11450
rect 11062 11398 11064 11450
rect 10902 11396 10926 11398
rect 10982 11396 11006 11398
rect 11062 11396 11086 11398
rect 10846 11376 11142 11396
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10612 5710 10640 11086
rect 11164 11082 11192 11154
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 9382 10732 10950
rect 10846 10364 11142 10384
rect 10902 10362 10926 10364
rect 10982 10362 11006 10364
rect 11062 10362 11086 10364
rect 10924 10310 10926 10362
rect 10988 10310 11000 10362
rect 11062 10310 11064 10362
rect 10902 10308 10926 10310
rect 10982 10308 11006 10310
rect 11062 10308 11086 10310
rect 10846 10288 11142 10308
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 10980 9722 11008 9998
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10846 9276 11142 9296
rect 10902 9274 10926 9276
rect 10982 9274 11006 9276
rect 11062 9274 11086 9276
rect 10924 9222 10926 9274
rect 10988 9222 11000 9274
rect 11062 9222 11064 9274
rect 10902 9220 10926 9222
rect 10982 9220 11006 9222
rect 11062 9220 11086 9222
rect 10846 9200 11142 9220
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10520 3466 10548 4082
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 10612 3126 10640 5238
rect 10704 3942 10732 8366
rect 10846 8188 11142 8208
rect 10902 8186 10926 8188
rect 10982 8186 11006 8188
rect 11062 8186 11086 8188
rect 10924 8134 10926 8186
rect 10988 8134 11000 8186
rect 11062 8134 11064 8186
rect 10902 8132 10926 8134
rect 10982 8132 11006 8134
rect 11062 8132 11086 8134
rect 10846 8112 11142 8132
rect 10846 7100 11142 7120
rect 10902 7098 10926 7100
rect 10982 7098 11006 7100
rect 11062 7098 11086 7100
rect 10924 7046 10926 7098
rect 10988 7046 11000 7098
rect 11062 7046 11064 7098
rect 10902 7044 10926 7046
rect 10982 7044 11006 7046
rect 11062 7044 11086 7046
rect 10846 7024 11142 7044
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6186 10824 6666
rect 11256 6254 11284 9318
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11244 6248 11296 6254
rect 11244 6190 11296 6196
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10846 6012 11142 6032
rect 10902 6010 10926 6012
rect 10982 6010 11006 6012
rect 11062 6010 11086 6012
rect 10924 5958 10926 6010
rect 10988 5958 11000 6010
rect 11062 5958 11064 6010
rect 10902 5956 10926 5958
rect 10982 5956 11006 5958
rect 11062 5956 11086 5958
rect 10846 5936 11142 5956
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10888 5710 10916 5743
rect 11256 5710 11284 6190
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10796 5545 10824 5578
rect 10782 5536 10838 5545
rect 10782 5471 10838 5480
rect 10888 5302 10916 5646
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 11256 5098 11284 5170
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 10846 4924 11142 4944
rect 10902 4922 10926 4924
rect 10982 4922 11006 4924
rect 11062 4922 11086 4924
rect 10924 4870 10926 4922
rect 10988 4870 11000 4922
rect 11062 4870 11064 4922
rect 10902 4868 10926 4870
rect 10982 4868 11006 4870
rect 11062 4868 11086 4870
rect 10846 4848 11142 4868
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10846 3836 11142 3856
rect 10902 3834 10926 3836
rect 10982 3834 11006 3836
rect 11062 3834 11086 3836
rect 10924 3782 10926 3834
rect 10988 3782 11000 3834
rect 11062 3782 11064 3834
rect 10902 3780 10926 3782
rect 10982 3780 11006 3782
rect 11062 3780 11086 3782
rect 10846 3760 11142 3780
rect 11348 3126 11376 9114
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11440 4622 11468 7346
rect 11532 6458 11560 9590
rect 11612 8832 11664 8838
rect 11612 8774 11664 8780
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11532 5681 11560 6190
rect 11518 5672 11574 5681
rect 11518 5607 11574 5616
rect 11624 4622 11652 8774
rect 11716 5914 11744 11698
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 10846 2748 11142 2768
rect 10902 2746 10926 2748
rect 10982 2746 11006 2748
rect 11062 2746 11086 2748
rect 10924 2694 10926 2746
rect 10988 2694 11000 2746
rect 11062 2694 11064 2746
rect 10902 2692 10926 2694
rect 10982 2692 11006 2694
rect 11062 2692 11086 2694
rect 10846 2672 11142 2692
rect 11440 2650 11468 4558
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11532 2582 11560 4490
rect 11624 2650 11652 4558
rect 11808 4078 11836 10610
rect 11900 10538 11928 12406
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 5624 11928 10474
rect 11992 7954 12020 12582
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11762 12112 12038
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12176 10266 12204 12702
rect 13464 12306 13492 15506
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 12254 11520 12310 11529
rect 12254 11455 12310 11464
rect 12268 11150 12296 11455
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 5778 12020 7890
rect 12176 6866 12204 10202
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12268 9625 12296 9998
rect 12254 9616 12310 9625
rect 12254 9551 12310 9560
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12268 7721 12296 7822
rect 12254 7712 12310 7721
rect 12254 7647 12310 7656
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12070 6760 12126 6769
rect 12070 6695 12072 6704
rect 12124 6695 12126 6704
rect 12072 6666 12124 6672
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 5817 12204 6598
rect 12162 5808 12218 5817
rect 11980 5772 12032 5778
rect 12162 5743 12218 5752
rect 11980 5714 12032 5720
rect 11980 5636 12032 5642
rect 11900 5596 11980 5624
rect 11980 5578 12032 5584
rect 11886 5400 11942 5409
rect 11886 5335 11942 5344
rect 11900 5302 11928 5335
rect 11888 5296 11940 5302
rect 11992 5273 12020 5578
rect 11888 5238 11940 5244
rect 11978 5264 12034 5273
rect 11978 5199 12034 5208
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4214 11928 4422
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11992 3602 12020 5034
rect 12162 3904 12218 3913
rect 12162 3839 12218 3848
rect 11980 3596 12032 3602
rect 11980 3538 12032 3544
rect 12176 3194 12204 3839
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 11520 2440 11572 2446
rect 11572 2400 11652 2428
rect 11520 2382 11572 2388
rect 10428 2009 10456 2382
rect 10414 2000 10470 2009
rect 10414 1935 10470 1944
rect 11624 800 11652 2400
rect 12912 800 12940 3470
rect 9678 96 9734 105
rect 9678 31 9734 40
rect 10322 0 10378 800
rect 11610 0 11666 800
rect 12898 0 12954 800
<< via2 >>
rect 1766 13388 1822 13424
rect 2778 15272 2834 15328
rect 1766 13368 1768 13388
rect 1768 13368 1820 13388
rect 1820 13368 1822 13388
rect 2934 13626 2990 13628
rect 3014 13626 3070 13628
rect 3094 13626 3150 13628
rect 3174 13626 3230 13628
rect 2934 13574 2960 13626
rect 2960 13574 2990 13626
rect 3014 13574 3024 13626
rect 3024 13574 3070 13626
rect 3094 13574 3140 13626
rect 3140 13574 3150 13626
rect 3174 13574 3204 13626
rect 3204 13574 3230 13626
rect 2934 13572 2990 13574
rect 3014 13572 3070 13574
rect 3094 13572 3150 13574
rect 3174 13572 3230 13574
rect 2934 12538 2990 12540
rect 3014 12538 3070 12540
rect 3094 12538 3150 12540
rect 3174 12538 3230 12540
rect 2934 12486 2960 12538
rect 2960 12486 2990 12538
rect 3014 12486 3024 12538
rect 3024 12486 3070 12538
rect 3094 12486 3140 12538
rect 3140 12486 3150 12538
rect 3174 12486 3204 12538
rect 3204 12486 3230 12538
rect 2934 12484 2990 12486
rect 3014 12484 3070 12486
rect 3094 12484 3150 12486
rect 3174 12484 3230 12486
rect 1398 11464 1454 11520
rect 1490 7692 1492 7712
rect 1492 7692 1544 7712
rect 1544 7692 1546 7712
rect 1490 7656 1546 7692
rect 1858 9560 1914 9616
rect 2934 11450 2990 11452
rect 3014 11450 3070 11452
rect 3094 11450 3150 11452
rect 3174 11450 3230 11452
rect 2934 11398 2960 11450
rect 2960 11398 2990 11450
rect 3014 11398 3024 11450
rect 3024 11398 3070 11450
rect 3094 11398 3140 11450
rect 3140 11398 3150 11450
rect 3174 11398 3204 11450
rect 3204 11398 3230 11450
rect 2934 11396 2990 11398
rect 3014 11396 3070 11398
rect 3094 11396 3150 11398
rect 3174 11396 3230 11398
rect 2934 10362 2990 10364
rect 3014 10362 3070 10364
rect 3094 10362 3150 10364
rect 3174 10362 3230 10364
rect 2934 10310 2960 10362
rect 2960 10310 2990 10362
rect 3014 10310 3024 10362
rect 3024 10310 3070 10362
rect 3094 10310 3140 10362
rect 3140 10310 3150 10362
rect 3174 10310 3204 10362
rect 3204 10310 3230 10362
rect 2934 10308 2990 10310
rect 3014 10308 3070 10310
rect 3094 10308 3150 10310
rect 3174 10308 3230 10310
rect 2934 9274 2990 9276
rect 3014 9274 3070 9276
rect 3094 9274 3150 9276
rect 3174 9274 3230 9276
rect 2934 9222 2960 9274
rect 2960 9222 2990 9274
rect 3014 9222 3024 9274
rect 3024 9222 3070 9274
rect 3094 9222 3140 9274
rect 3140 9222 3150 9274
rect 3174 9222 3204 9274
rect 3204 9222 3230 9274
rect 2934 9220 2990 9222
rect 3014 9220 3070 9222
rect 3094 9220 3150 9222
rect 3174 9220 3230 9222
rect 2934 8186 2990 8188
rect 3014 8186 3070 8188
rect 3094 8186 3150 8188
rect 3174 8186 3230 8188
rect 2934 8134 2960 8186
rect 2960 8134 2990 8186
rect 3014 8134 3024 8186
rect 3024 8134 3070 8186
rect 3094 8134 3140 8186
rect 3140 8134 3150 8186
rect 3174 8134 3204 8186
rect 3204 8134 3230 8186
rect 2934 8132 2990 8134
rect 3014 8132 3070 8134
rect 3094 8132 3150 8134
rect 3174 8132 3230 8134
rect 1398 5752 1454 5808
rect 2410 6704 2466 6760
rect 2934 7098 2990 7100
rect 3014 7098 3070 7100
rect 3094 7098 3150 7100
rect 3174 7098 3230 7100
rect 2934 7046 2960 7098
rect 2960 7046 2990 7098
rect 3014 7046 3024 7098
rect 3024 7046 3070 7098
rect 3094 7046 3140 7098
rect 3140 7046 3150 7098
rect 3174 7046 3204 7098
rect 3204 7046 3230 7098
rect 2934 7044 2990 7046
rect 3014 7044 3070 7046
rect 3094 7044 3150 7046
rect 3174 7044 3230 7046
rect 2934 6010 2990 6012
rect 3014 6010 3070 6012
rect 3094 6010 3150 6012
rect 3174 6010 3230 6012
rect 2934 5958 2960 6010
rect 2960 5958 2990 6010
rect 3014 5958 3024 6010
rect 3024 5958 3070 6010
rect 3094 5958 3140 6010
rect 3140 5958 3150 6010
rect 3174 5958 3204 6010
rect 3204 5958 3230 6010
rect 2934 5956 2990 5958
rect 3014 5956 3070 5958
rect 3094 5956 3150 5958
rect 3174 5956 3230 5958
rect 2934 4922 2990 4924
rect 3014 4922 3070 4924
rect 3094 4922 3150 4924
rect 3174 4922 3230 4924
rect 2934 4870 2960 4922
rect 2960 4870 2990 4922
rect 3014 4870 3024 4922
rect 3024 4870 3070 4922
rect 3094 4870 3140 4922
rect 3140 4870 3150 4922
rect 3174 4870 3204 4922
rect 3204 4870 3230 4922
rect 2934 4868 2990 4870
rect 3014 4868 3070 4870
rect 3094 4868 3150 4870
rect 3174 4868 3230 4870
rect 1858 3884 1860 3904
rect 1860 3884 1912 3904
rect 1912 3884 1914 3904
rect 1858 3848 1914 3884
rect 2934 3834 2990 3836
rect 3014 3834 3070 3836
rect 3094 3834 3150 3836
rect 3174 3834 3230 3836
rect 2934 3782 2960 3834
rect 2960 3782 2990 3834
rect 3014 3782 3024 3834
rect 3024 3782 3070 3834
rect 3094 3782 3140 3834
rect 3140 3782 3150 3834
rect 3174 3782 3204 3834
rect 3204 3782 3230 3834
rect 2934 3780 2990 3782
rect 3014 3780 3070 3782
rect 3094 3780 3150 3782
rect 3174 3780 3230 3782
rect 3790 12180 3792 12200
rect 3792 12180 3844 12200
rect 3844 12180 3846 12200
rect 3790 12144 3846 12180
rect 4342 12180 4344 12200
rect 4344 12180 4396 12200
rect 4396 12180 4398 12200
rect 4342 12144 4398 12180
rect 4912 13082 4968 13084
rect 4992 13082 5048 13084
rect 5072 13082 5128 13084
rect 5152 13082 5208 13084
rect 4912 13030 4938 13082
rect 4938 13030 4968 13082
rect 4992 13030 5002 13082
rect 5002 13030 5048 13082
rect 5072 13030 5118 13082
rect 5118 13030 5128 13082
rect 5152 13030 5182 13082
rect 5182 13030 5208 13082
rect 4912 13028 4968 13030
rect 4992 13028 5048 13030
rect 5072 13028 5128 13030
rect 5152 13028 5208 13030
rect 4434 6296 4490 6352
rect 4434 6160 4490 6216
rect 4710 11600 4766 11656
rect 4912 11994 4968 11996
rect 4992 11994 5048 11996
rect 5072 11994 5128 11996
rect 5152 11994 5208 11996
rect 4912 11942 4938 11994
rect 4938 11942 4968 11994
rect 4992 11942 5002 11994
rect 5002 11942 5048 11994
rect 5072 11942 5118 11994
rect 5118 11942 5128 11994
rect 5152 11942 5182 11994
rect 5182 11942 5208 11994
rect 4912 11940 4968 11942
rect 4992 11940 5048 11942
rect 5072 11940 5128 11942
rect 5152 11940 5208 11942
rect 4912 10906 4968 10908
rect 4992 10906 5048 10908
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 4912 10854 4938 10906
rect 4938 10854 4968 10906
rect 4992 10854 5002 10906
rect 5002 10854 5048 10906
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5208 10906
rect 4912 10852 4968 10854
rect 4992 10852 5048 10854
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 4912 9818 4968 9820
rect 4992 9818 5048 9820
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 4912 9766 4938 9818
rect 4938 9766 4968 9818
rect 4992 9766 5002 9818
rect 5002 9766 5048 9818
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5208 9818
rect 4912 9764 4968 9766
rect 4992 9764 5048 9766
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 4912 8730 4968 8732
rect 4992 8730 5048 8732
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 4912 8678 4938 8730
rect 4938 8678 4968 8730
rect 4992 8678 5002 8730
rect 5002 8678 5048 8730
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5208 8730
rect 4912 8676 4968 8678
rect 4992 8676 5048 8678
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 4912 7642 4968 7644
rect 4992 7642 5048 7644
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 4912 7590 4938 7642
rect 4938 7590 4968 7642
rect 4992 7590 5002 7642
rect 5002 7590 5048 7642
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5208 7642
rect 4912 7588 4968 7590
rect 4992 7588 5048 7590
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 4912 6554 4968 6556
rect 4992 6554 5048 6556
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 4912 6502 4938 6554
rect 4938 6502 4968 6554
rect 4992 6502 5002 6554
rect 5002 6502 5048 6554
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5208 6554
rect 4912 6500 4968 6502
rect 4992 6500 5048 6502
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 4912 5466 4968 5468
rect 4992 5466 5048 5468
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 4912 5414 4938 5466
rect 4938 5414 4968 5466
rect 4992 5414 5002 5466
rect 5002 5414 5048 5466
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5208 5466
rect 4912 5412 4968 5414
rect 4992 5412 5048 5414
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 6890 13626 6946 13628
rect 6970 13626 7026 13628
rect 7050 13626 7106 13628
rect 7130 13626 7186 13628
rect 6890 13574 6916 13626
rect 6916 13574 6946 13626
rect 6970 13574 6980 13626
rect 6980 13574 7026 13626
rect 7050 13574 7096 13626
rect 7096 13574 7106 13626
rect 7130 13574 7160 13626
rect 7160 13574 7186 13626
rect 6890 13572 6946 13574
rect 6970 13572 7026 13574
rect 7050 13572 7106 13574
rect 7130 13572 7186 13574
rect 6890 12538 6946 12540
rect 6970 12538 7026 12540
rect 7050 12538 7106 12540
rect 7130 12538 7186 12540
rect 6890 12486 6916 12538
rect 6916 12486 6946 12538
rect 6970 12486 6980 12538
rect 6980 12486 7026 12538
rect 7050 12486 7096 12538
rect 7096 12486 7106 12538
rect 7130 12486 7160 12538
rect 7160 12486 7186 12538
rect 6890 12484 6946 12486
rect 6970 12484 7026 12486
rect 7050 12484 7106 12486
rect 7130 12484 7186 12486
rect 4912 4378 4968 4380
rect 4992 4378 5048 4380
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 4912 4326 4938 4378
rect 4938 4326 4968 4378
rect 4992 4326 5002 4378
rect 5002 4326 5048 4378
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5208 4378
rect 4912 4324 4968 4326
rect 4992 4324 5048 4326
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 4912 3290 4968 3292
rect 4992 3290 5048 3292
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 4912 3238 4938 3290
rect 4938 3238 4968 3290
rect 4992 3238 5002 3290
rect 5002 3238 5048 3290
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5208 3290
rect 4912 3236 4968 3238
rect 4992 3236 5048 3238
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 2934 2746 2990 2748
rect 3014 2746 3070 2748
rect 3094 2746 3150 2748
rect 3174 2746 3230 2748
rect 2934 2694 2960 2746
rect 2960 2694 2990 2746
rect 3014 2694 3024 2746
rect 3024 2694 3070 2746
rect 3094 2694 3140 2746
rect 3140 2694 3150 2746
rect 3174 2694 3204 2746
rect 3204 2694 3230 2746
rect 2934 2692 2990 2694
rect 3014 2692 3070 2694
rect 3094 2692 3150 2694
rect 3174 2692 3230 2694
rect 5814 5228 5870 5264
rect 5814 5208 5816 5228
rect 5816 5208 5868 5228
rect 5868 5208 5870 5228
rect 6918 11600 6974 11656
rect 6890 11450 6946 11452
rect 6970 11450 7026 11452
rect 7050 11450 7106 11452
rect 7130 11450 7186 11452
rect 6890 11398 6916 11450
rect 6916 11398 6946 11450
rect 6970 11398 6980 11450
rect 6980 11398 7026 11450
rect 7050 11398 7096 11450
rect 7096 11398 7106 11450
rect 7130 11398 7160 11450
rect 7160 11398 7186 11450
rect 6890 11396 6946 11398
rect 6970 11396 7026 11398
rect 7050 11396 7106 11398
rect 7130 11396 7186 11398
rect 6890 10362 6946 10364
rect 6970 10362 7026 10364
rect 7050 10362 7106 10364
rect 7130 10362 7186 10364
rect 6890 10310 6916 10362
rect 6916 10310 6946 10362
rect 6970 10310 6980 10362
rect 6980 10310 7026 10362
rect 7050 10310 7096 10362
rect 7096 10310 7106 10362
rect 7130 10310 7160 10362
rect 7160 10310 7186 10362
rect 6890 10308 6946 10310
rect 6970 10308 7026 10310
rect 7050 10308 7106 10310
rect 7130 10308 7186 10310
rect 6890 9274 6946 9276
rect 6970 9274 7026 9276
rect 7050 9274 7106 9276
rect 7130 9274 7186 9276
rect 6890 9222 6916 9274
rect 6916 9222 6946 9274
rect 6970 9222 6980 9274
rect 6980 9222 7026 9274
rect 7050 9222 7096 9274
rect 7096 9222 7106 9274
rect 7130 9222 7160 9274
rect 7160 9222 7186 9274
rect 6890 9220 6946 9222
rect 6970 9220 7026 9222
rect 7050 9220 7106 9222
rect 7130 9220 7186 9222
rect 6890 8186 6946 8188
rect 6970 8186 7026 8188
rect 7050 8186 7106 8188
rect 7130 8186 7186 8188
rect 6890 8134 6916 8186
rect 6916 8134 6946 8186
rect 6970 8134 6980 8186
rect 6980 8134 7026 8186
rect 7050 8134 7096 8186
rect 7096 8134 7106 8186
rect 7130 8134 7160 8186
rect 7160 8134 7186 8186
rect 6890 8132 6946 8134
rect 6970 8132 7026 8134
rect 7050 8132 7106 8134
rect 7130 8132 7186 8134
rect 8868 13082 8924 13084
rect 8948 13082 9004 13084
rect 9028 13082 9084 13084
rect 9108 13082 9164 13084
rect 8868 13030 8894 13082
rect 8894 13030 8924 13082
rect 8948 13030 8958 13082
rect 8958 13030 9004 13082
rect 9028 13030 9074 13082
rect 9074 13030 9084 13082
rect 9108 13030 9138 13082
rect 9138 13030 9164 13082
rect 8868 13028 8924 13030
rect 8948 13028 9004 13030
rect 9028 13028 9084 13030
rect 9108 13028 9164 13030
rect 6890 7098 6946 7100
rect 6970 7098 7026 7100
rect 7050 7098 7106 7100
rect 7130 7098 7186 7100
rect 6890 7046 6916 7098
rect 6916 7046 6946 7098
rect 6970 7046 6980 7098
rect 6980 7046 7026 7098
rect 7050 7046 7096 7098
rect 7096 7046 7106 7098
rect 7130 7046 7160 7098
rect 7160 7046 7186 7098
rect 6890 7044 6946 7046
rect 6970 7044 7026 7046
rect 7050 7044 7106 7046
rect 7130 7044 7186 7046
rect 6734 6296 6790 6352
rect 7102 6840 7158 6896
rect 7194 6432 7250 6488
rect 6890 6010 6946 6012
rect 6970 6010 7026 6012
rect 7050 6010 7106 6012
rect 7130 6010 7186 6012
rect 6890 5958 6916 6010
rect 6916 5958 6946 6010
rect 6970 5958 6980 6010
rect 6980 5958 7026 6010
rect 7050 5958 7096 6010
rect 7096 5958 7106 6010
rect 7130 5958 7160 6010
rect 7160 5958 7186 6010
rect 6890 5956 6946 5958
rect 6970 5956 7026 5958
rect 7050 5956 7106 5958
rect 7130 5956 7186 5958
rect 6826 5772 6882 5808
rect 6826 5752 6828 5772
rect 6828 5752 6880 5772
rect 6880 5752 6882 5772
rect 6890 4922 6946 4924
rect 6970 4922 7026 4924
rect 7050 4922 7106 4924
rect 7130 4922 7186 4924
rect 6890 4870 6916 4922
rect 6916 4870 6946 4922
rect 6970 4870 6980 4922
rect 6980 4870 7026 4922
rect 7050 4870 7096 4922
rect 7096 4870 7106 4922
rect 7130 4870 7160 4922
rect 7160 4870 7186 4922
rect 6890 4868 6946 4870
rect 6970 4868 7026 4870
rect 7050 4868 7106 4870
rect 7130 4868 7186 4870
rect 6890 3834 6946 3836
rect 6970 3834 7026 3836
rect 7050 3834 7106 3836
rect 7130 3834 7186 3836
rect 6890 3782 6916 3834
rect 6916 3782 6946 3834
rect 6970 3782 6980 3834
rect 6980 3782 7026 3834
rect 7050 3782 7096 3834
rect 7096 3782 7106 3834
rect 7130 3782 7160 3834
rect 7160 3782 7186 3834
rect 6890 3780 6946 3782
rect 6970 3780 7026 3782
rect 7050 3780 7106 3782
rect 7130 3780 7186 3782
rect 6890 2746 6946 2748
rect 6970 2746 7026 2748
rect 7050 2746 7106 2748
rect 7130 2746 7186 2748
rect 6890 2694 6916 2746
rect 6916 2694 6946 2746
rect 6970 2694 6980 2746
rect 6980 2694 7026 2746
rect 7050 2694 7096 2746
rect 7096 2694 7106 2746
rect 7130 2694 7160 2746
rect 7160 2694 7186 2746
rect 6890 2692 6946 2694
rect 6970 2692 7026 2694
rect 7050 2692 7106 2694
rect 7130 2692 7186 2694
rect 10598 15272 10654 15328
rect 8868 11994 8924 11996
rect 8948 11994 9004 11996
rect 9028 11994 9084 11996
rect 9108 11994 9164 11996
rect 8868 11942 8894 11994
rect 8894 11942 8924 11994
rect 8948 11942 8958 11994
rect 8958 11942 9004 11994
rect 9028 11942 9074 11994
rect 9074 11942 9084 11994
rect 9108 11942 9138 11994
rect 9138 11942 9164 11994
rect 8868 11940 8924 11942
rect 8948 11940 9004 11942
rect 9028 11940 9084 11942
rect 9108 11940 9164 11942
rect 7746 7112 7802 7168
rect 7562 5616 7618 5672
rect 1398 1944 1454 2000
rect 4912 2202 4968 2204
rect 4992 2202 5048 2204
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 4912 2150 4938 2202
rect 4938 2150 4968 2202
rect 4992 2150 5002 2202
rect 5002 2150 5048 2202
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5208 2202
rect 4912 2148 4968 2150
rect 4992 2148 5048 2150
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 8868 10906 8924 10908
rect 8948 10906 9004 10908
rect 9028 10906 9084 10908
rect 9108 10906 9164 10908
rect 8868 10854 8894 10906
rect 8894 10854 8924 10906
rect 8948 10854 8958 10906
rect 8958 10854 9004 10906
rect 9028 10854 9074 10906
rect 9074 10854 9084 10906
rect 9108 10854 9138 10906
rect 9138 10854 9164 10906
rect 8868 10852 8924 10854
rect 8948 10852 9004 10854
rect 9028 10852 9084 10854
rect 9108 10852 9164 10854
rect 8574 6432 8630 6488
rect 8868 9818 8924 9820
rect 8948 9818 9004 9820
rect 9028 9818 9084 9820
rect 9108 9818 9164 9820
rect 8868 9766 8894 9818
rect 8894 9766 8924 9818
rect 8948 9766 8958 9818
rect 8958 9766 9004 9818
rect 9028 9766 9074 9818
rect 9074 9766 9084 9818
rect 9108 9766 9138 9818
rect 9138 9766 9164 9818
rect 8868 9764 8924 9766
rect 8948 9764 9004 9766
rect 9028 9764 9084 9766
rect 9108 9764 9164 9766
rect 8868 8730 8924 8732
rect 8948 8730 9004 8732
rect 9028 8730 9084 8732
rect 9108 8730 9164 8732
rect 8868 8678 8894 8730
rect 8894 8678 8924 8730
rect 8948 8678 8958 8730
rect 8958 8678 9004 8730
rect 9028 8678 9074 8730
rect 9074 8678 9084 8730
rect 9108 8678 9138 8730
rect 9138 8678 9164 8730
rect 8868 8676 8924 8678
rect 8948 8676 9004 8678
rect 9028 8676 9084 8678
rect 9108 8676 9164 8678
rect 8868 7642 8924 7644
rect 8948 7642 9004 7644
rect 9028 7642 9084 7644
rect 9108 7642 9164 7644
rect 8868 7590 8894 7642
rect 8894 7590 8924 7642
rect 8948 7590 8958 7642
rect 8958 7590 9004 7642
rect 9028 7590 9074 7642
rect 9074 7590 9084 7642
rect 9108 7590 9138 7642
rect 9138 7590 9164 7642
rect 8868 7588 8924 7590
rect 8948 7588 9004 7590
rect 9028 7588 9084 7590
rect 9108 7588 9164 7590
rect 8850 6840 8906 6896
rect 8868 6554 8924 6556
rect 8948 6554 9004 6556
rect 9028 6554 9084 6556
rect 9108 6554 9164 6556
rect 8868 6502 8894 6554
rect 8894 6502 8924 6554
rect 8948 6502 8958 6554
rect 8958 6502 9004 6554
rect 9028 6502 9074 6554
rect 9074 6502 9084 6554
rect 9108 6502 9138 6554
rect 9138 6502 9164 6554
rect 8868 6500 8924 6502
rect 8948 6500 9004 6502
rect 9028 6500 9084 6502
rect 9108 6500 9164 6502
rect 9034 6180 9090 6216
rect 9034 6160 9036 6180
rect 9036 6160 9088 6180
rect 9088 6160 9090 6180
rect 8868 5466 8924 5468
rect 8948 5466 9004 5468
rect 9028 5466 9084 5468
rect 9108 5466 9164 5468
rect 8868 5414 8894 5466
rect 8894 5414 8924 5466
rect 8948 5414 8958 5466
rect 8958 5414 9004 5466
rect 9028 5414 9074 5466
rect 9074 5414 9084 5466
rect 9108 5414 9138 5466
rect 9138 5414 9164 5466
rect 8868 5412 8924 5414
rect 8948 5412 9004 5414
rect 9028 5412 9084 5414
rect 9108 5412 9164 5414
rect 8868 4378 8924 4380
rect 8948 4378 9004 4380
rect 9028 4378 9084 4380
rect 9108 4378 9164 4380
rect 8868 4326 8894 4378
rect 8894 4326 8924 4378
rect 8948 4326 8958 4378
rect 8958 4326 9004 4378
rect 9028 4326 9074 4378
rect 9074 4326 9084 4378
rect 9108 4326 9138 4378
rect 9138 4326 9164 4378
rect 8868 4324 8924 4326
rect 8948 4324 9004 4326
rect 9028 4324 9084 4326
rect 9108 4324 9164 4326
rect 8868 3290 8924 3292
rect 8948 3290 9004 3292
rect 9028 3290 9084 3292
rect 9108 3290 9164 3292
rect 8868 3238 8894 3290
rect 8894 3238 8924 3290
rect 8948 3238 8958 3290
rect 8958 3238 9004 3290
rect 9028 3238 9074 3290
rect 9074 3238 9084 3290
rect 9108 3238 9138 3290
rect 9138 3238 9164 3290
rect 8868 3236 8924 3238
rect 8948 3236 9004 3238
rect 9028 3236 9084 3238
rect 9108 3236 9164 3238
rect 9678 6568 9734 6624
rect 9862 6568 9918 6624
rect 9954 6432 10010 6488
rect 9954 6296 10010 6352
rect 9862 6160 9918 6216
rect 9678 5888 9734 5944
rect 9586 5208 9642 5264
rect 8868 2202 8924 2204
rect 8948 2202 9004 2204
rect 9028 2202 9084 2204
rect 9108 2202 9164 2204
rect 8868 2150 8894 2202
rect 8894 2150 8924 2202
rect 8948 2150 8958 2202
rect 8958 2150 9004 2202
rect 9028 2150 9074 2202
rect 9074 2150 9084 2202
rect 9108 2150 9138 2202
rect 9138 2150 9164 2202
rect 8868 2148 8924 2150
rect 8948 2148 9004 2150
rect 9028 2148 9084 2150
rect 9108 2148 9164 2150
rect 9770 5344 9826 5400
rect 10230 5480 10286 5536
rect 10138 5208 10194 5264
rect 10414 6316 10470 6352
rect 10414 6296 10416 6316
rect 10416 6296 10468 6316
rect 10468 6296 10470 6316
rect 9954 4004 10010 4040
rect 9954 3984 9956 4004
rect 9956 3984 10008 4004
rect 10008 3984 10010 4004
rect 10846 13626 10902 13628
rect 10926 13626 10982 13628
rect 11006 13626 11062 13628
rect 11086 13626 11142 13628
rect 10846 13574 10872 13626
rect 10872 13574 10902 13626
rect 10926 13574 10936 13626
rect 10936 13574 10982 13626
rect 11006 13574 11052 13626
rect 11052 13574 11062 13626
rect 11086 13574 11116 13626
rect 11116 13574 11142 13626
rect 10846 13572 10902 13574
rect 10926 13572 10982 13574
rect 11006 13572 11062 13574
rect 11086 13572 11142 13574
rect 10966 13388 11022 13424
rect 10966 13368 10968 13388
rect 10968 13368 11020 13388
rect 11020 13368 11022 13388
rect 10846 12538 10902 12540
rect 10926 12538 10982 12540
rect 11006 12538 11062 12540
rect 11086 12538 11142 12540
rect 10846 12486 10872 12538
rect 10872 12486 10902 12538
rect 10926 12486 10936 12538
rect 10936 12486 10982 12538
rect 11006 12486 11052 12538
rect 11052 12486 11062 12538
rect 11086 12486 11116 12538
rect 11116 12486 11142 12538
rect 10846 12484 10902 12486
rect 10926 12484 10982 12486
rect 11006 12484 11062 12486
rect 11086 12484 11142 12486
rect 10846 11450 10902 11452
rect 10926 11450 10982 11452
rect 11006 11450 11062 11452
rect 11086 11450 11142 11452
rect 10846 11398 10872 11450
rect 10872 11398 10902 11450
rect 10926 11398 10936 11450
rect 10936 11398 10982 11450
rect 11006 11398 11052 11450
rect 11052 11398 11062 11450
rect 11086 11398 11116 11450
rect 11116 11398 11142 11450
rect 10846 11396 10902 11398
rect 10926 11396 10982 11398
rect 11006 11396 11062 11398
rect 11086 11396 11142 11398
rect 10846 10362 10902 10364
rect 10926 10362 10982 10364
rect 11006 10362 11062 10364
rect 11086 10362 11142 10364
rect 10846 10310 10872 10362
rect 10872 10310 10902 10362
rect 10926 10310 10936 10362
rect 10936 10310 10982 10362
rect 11006 10310 11052 10362
rect 11052 10310 11062 10362
rect 11086 10310 11116 10362
rect 11116 10310 11142 10362
rect 10846 10308 10902 10310
rect 10926 10308 10982 10310
rect 11006 10308 11062 10310
rect 11086 10308 11142 10310
rect 10846 9274 10902 9276
rect 10926 9274 10982 9276
rect 11006 9274 11062 9276
rect 11086 9274 11142 9276
rect 10846 9222 10872 9274
rect 10872 9222 10902 9274
rect 10926 9222 10936 9274
rect 10936 9222 10982 9274
rect 11006 9222 11052 9274
rect 11052 9222 11062 9274
rect 11086 9222 11116 9274
rect 11116 9222 11142 9274
rect 10846 9220 10902 9222
rect 10926 9220 10982 9222
rect 11006 9220 11062 9222
rect 11086 9220 11142 9222
rect 10846 8186 10902 8188
rect 10926 8186 10982 8188
rect 11006 8186 11062 8188
rect 11086 8186 11142 8188
rect 10846 8134 10872 8186
rect 10872 8134 10902 8186
rect 10926 8134 10936 8186
rect 10936 8134 10982 8186
rect 11006 8134 11052 8186
rect 11052 8134 11062 8186
rect 11086 8134 11116 8186
rect 11116 8134 11142 8186
rect 10846 8132 10902 8134
rect 10926 8132 10982 8134
rect 11006 8132 11062 8134
rect 11086 8132 11142 8134
rect 10846 7098 10902 7100
rect 10926 7098 10982 7100
rect 11006 7098 11062 7100
rect 11086 7098 11142 7100
rect 10846 7046 10872 7098
rect 10872 7046 10902 7098
rect 10926 7046 10936 7098
rect 10936 7046 10982 7098
rect 11006 7046 11052 7098
rect 11052 7046 11062 7098
rect 11086 7046 11116 7098
rect 11116 7046 11142 7098
rect 10846 7044 10902 7046
rect 10926 7044 10982 7046
rect 11006 7044 11062 7046
rect 11086 7044 11142 7046
rect 10846 6010 10902 6012
rect 10926 6010 10982 6012
rect 11006 6010 11062 6012
rect 11086 6010 11142 6012
rect 10846 5958 10872 6010
rect 10872 5958 10902 6010
rect 10926 5958 10936 6010
rect 10936 5958 10982 6010
rect 11006 5958 11052 6010
rect 11052 5958 11062 6010
rect 11086 5958 11116 6010
rect 11116 5958 11142 6010
rect 10846 5956 10902 5958
rect 10926 5956 10982 5958
rect 11006 5956 11062 5958
rect 11086 5956 11142 5958
rect 10874 5752 10930 5808
rect 10782 5480 10838 5536
rect 10846 4922 10902 4924
rect 10926 4922 10982 4924
rect 11006 4922 11062 4924
rect 11086 4922 11142 4924
rect 10846 4870 10872 4922
rect 10872 4870 10902 4922
rect 10926 4870 10936 4922
rect 10936 4870 10982 4922
rect 11006 4870 11052 4922
rect 11052 4870 11062 4922
rect 11086 4870 11116 4922
rect 11116 4870 11142 4922
rect 10846 4868 10902 4870
rect 10926 4868 10982 4870
rect 11006 4868 11062 4870
rect 11086 4868 11142 4870
rect 10846 3834 10902 3836
rect 10926 3834 10982 3836
rect 11006 3834 11062 3836
rect 11086 3834 11142 3836
rect 10846 3782 10872 3834
rect 10872 3782 10902 3834
rect 10926 3782 10936 3834
rect 10936 3782 10982 3834
rect 11006 3782 11052 3834
rect 11052 3782 11062 3834
rect 11086 3782 11116 3834
rect 11116 3782 11142 3834
rect 10846 3780 10902 3782
rect 10926 3780 10982 3782
rect 11006 3780 11062 3782
rect 11086 3780 11142 3782
rect 11518 5616 11574 5672
rect 10846 2746 10902 2748
rect 10926 2746 10982 2748
rect 11006 2746 11062 2748
rect 11086 2746 11142 2748
rect 10846 2694 10872 2746
rect 10872 2694 10902 2746
rect 10926 2694 10936 2746
rect 10936 2694 10982 2746
rect 11006 2694 11052 2746
rect 11052 2694 11062 2746
rect 11086 2694 11116 2746
rect 11116 2694 11142 2746
rect 10846 2692 10902 2694
rect 10926 2692 10982 2694
rect 11006 2692 11062 2694
rect 11086 2692 11142 2694
rect 12254 11464 12310 11520
rect 12254 9560 12310 9616
rect 12254 7656 12310 7712
rect 12070 6724 12126 6760
rect 12070 6704 12072 6724
rect 12072 6704 12124 6724
rect 12124 6704 12126 6724
rect 12162 5752 12218 5808
rect 11886 5344 11942 5400
rect 11978 5208 12034 5264
rect 12162 3848 12218 3904
rect 10414 1944 10470 2000
rect 9678 40 9734 96
<< metal3 >>
rect 0 15330 800 15360
rect 2773 15330 2839 15333
rect 0 15328 2839 15330
rect 0 15272 2778 15328
rect 2834 15272 2839 15328
rect 0 15270 2839 15272
rect 0 15240 800 15270
rect 2773 15267 2839 15270
rect 10593 15330 10659 15333
rect 13362 15330 14162 15360
rect 10593 15328 14162 15330
rect 10593 15272 10598 15328
rect 10654 15272 14162 15328
rect 10593 15270 14162 15272
rect 10593 15267 10659 15270
rect 13362 15240 14162 15270
rect 2922 13632 3242 13633
rect 2922 13568 2930 13632
rect 2994 13568 3010 13632
rect 3074 13568 3090 13632
rect 3154 13568 3170 13632
rect 3234 13568 3242 13632
rect 2922 13567 3242 13568
rect 6878 13632 7198 13633
rect 6878 13568 6886 13632
rect 6950 13568 6966 13632
rect 7030 13568 7046 13632
rect 7110 13568 7126 13632
rect 7190 13568 7198 13632
rect 6878 13567 7198 13568
rect 10834 13632 11154 13633
rect 10834 13568 10842 13632
rect 10906 13568 10922 13632
rect 10986 13568 11002 13632
rect 11066 13568 11082 13632
rect 11146 13568 11154 13632
rect 10834 13567 11154 13568
rect 0 13426 800 13456
rect 1761 13426 1827 13429
rect 0 13424 1827 13426
rect 0 13368 1766 13424
rect 1822 13368 1827 13424
rect 0 13366 1827 13368
rect 0 13336 800 13366
rect 1761 13363 1827 13366
rect 10961 13426 11027 13429
rect 13362 13426 14162 13456
rect 10961 13424 14162 13426
rect 10961 13368 10966 13424
rect 11022 13368 14162 13424
rect 10961 13366 14162 13368
rect 10961 13363 11027 13366
rect 13362 13336 14162 13366
rect 4900 13088 5220 13089
rect 4900 13024 4908 13088
rect 4972 13024 4988 13088
rect 5052 13024 5068 13088
rect 5132 13024 5148 13088
rect 5212 13024 5220 13088
rect 4900 13023 5220 13024
rect 8856 13088 9176 13089
rect 8856 13024 8864 13088
rect 8928 13024 8944 13088
rect 9008 13024 9024 13088
rect 9088 13024 9104 13088
rect 9168 13024 9176 13088
rect 8856 13023 9176 13024
rect 2922 12544 3242 12545
rect 2922 12480 2930 12544
rect 2994 12480 3010 12544
rect 3074 12480 3090 12544
rect 3154 12480 3170 12544
rect 3234 12480 3242 12544
rect 2922 12479 3242 12480
rect 6878 12544 7198 12545
rect 6878 12480 6886 12544
rect 6950 12480 6966 12544
rect 7030 12480 7046 12544
rect 7110 12480 7126 12544
rect 7190 12480 7198 12544
rect 6878 12479 7198 12480
rect 10834 12544 11154 12545
rect 10834 12480 10842 12544
rect 10906 12480 10922 12544
rect 10986 12480 11002 12544
rect 11066 12480 11082 12544
rect 11146 12480 11154 12544
rect 10834 12479 11154 12480
rect 3785 12202 3851 12205
rect 4337 12202 4403 12205
rect 3785 12200 4403 12202
rect 3785 12144 3790 12200
rect 3846 12144 4342 12200
rect 4398 12144 4403 12200
rect 3785 12142 4403 12144
rect 3785 12139 3851 12142
rect 4337 12139 4403 12142
rect 4900 12000 5220 12001
rect 4900 11936 4908 12000
rect 4972 11936 4988 12000
rect 5052 11936 5068 12000
rect 5132 11936 5148 12000
rect 5212 11936 5220 12000
rect 4900 11935 5220 11936
rect 8856 12000 9176 12001
rect 8856 11936 8864 12000
rect 8928 11936 8944 12000
rect 9008 11936 9024 12000
rect 9088 11936 9104 12000
rect 9168 11936 9176 12000
rect 8856 11935 9176 11936
rect 4705 11658 4771 11661
rect 6913 11658 6979 11661
rect 4705 11656 6979 11658
rect 4705 11600 4710 11656
rect 4766 11600 6918 11656
rect 6974 11600 6979 11656
rect 4705 11598 6979 11600
rect 4705 11595 4771 11598
rect 6913 11595 6979 11598
rect 0 11522 800 11552
rect 1393 11522 1459 11525
rect 0 11520 1459 11522
rect 0 11464 1398 11520
rect 1454 11464 1459 11520
rect 0 11462 1459 11464
rect 0 11432 800 11462
rect 1393 11459 1459 11462
rect 12249 11522 12315 11525
rect 13362 11522 14162 11552
rect 12249 11520 14162 11522
rect 12249 11464 12254 11520
rect 12310 11464 14162 11520
rect 12249 11462 14162 11464
rect 12249 11459 12315 11462
rect 2922 11456 3242 11457
rect 2922 11392 2930 11456
rect 2994 11392 3010 11456
rect 3074 11392 3090 11456
rect 3154 11392 3170 11456
rect 3234 11392 3242 11456
rect 2922 11391 3242 11392
rect 6878 11456 7198 11457
rect 6878 11392 6886 11456
rect 6950 11392 6966 11456
rect 7030 11392 7046 11456
rect 7110 11392 7126 11456
rect 7190 11392 7198 11456
rect 6878 11391 7198 11392
rect 10834 11456 11154 11457
rect 10834 11392 10842 11456
rect 10906 11392 10922 11456
rect 10986 11392 11002 11456
rect 11066 11392 11082 11456
rect 11146 11392 11154 11456
rect 13362 11432 14162 11462
rect 10834 11391 11154 11392
rect 4900 10912 5220 10913
rect 4900 10848 4908 10912
rect 4972 10848 4988 10912
rect 5052 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5220 10912
rect 4900 10847 5220 10848
rect 8856 10912 9176 10913
rect 8856 10848 8864 10912
rect 8928 10848 8944 10912
rect 9008 10848 9024 10912
rect 9088 10848 9104 10912
rect 9168 10848 9176 10912
rect 8856 10847 9176 10848
rect 2922 10368 3242 10369
rect 2922 10304 2930 10368
rect 2994 10304 3010 10368
rect 3074 10304 3090 10368
rect 3154 10304 3170 10368
rect 3234 10304 3242 10368
rect 2922 10303 3242 10304
rect 6878 10368 7198 10369
rect 6878 10304 6886 10368
rect 6950 10304 6966 10368
rect 7030 10304 7046 10368
rect 7110 10304 7126 10368
rect 7190 10304 7198 10368
rect 6878 10303 7198 10304
rect 10834 10368 11154 10369
rect 10834 10304 10842 10368
rect 10906 10304 10922 10368
rect 10986 10304 11002 10368
rect 11066 10304 11082 10368
rect 11146 10304 11154 10368
rect 10834 10303 11154 10304
rect 4900 9824 5220 9825
rect 4900 9760 4908 9824
rect 4972 9760 4988 9824
rect 5052 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5220 9824
rect 4900 9759 5220 9760
rect 8856 9824 9176 9825
rect 8856 9760 8864 9824
rect 8928 9760 8944 9824
rect 9008 9760 9024 9824
rect 9088 9760 9104 9824
rect 9168 9760 9176 9824
rect 8856 9759 9176 9760
rect 0 9618 800 9648
rect 1853 9618 1919 9621
rect 0 9616 1919 9618
rect 0 9560 1858 9616
rect 1914 9560 1919 9616
rect 0 9558 1919 9560
rect 0 9528 800 9558
rect 1853 9555 1919 9558
rect 12249 9618 12315 9621
rect 13362 9618 14162 9648
rect 12249 9616 14162 9618
rect 12249 9560 12254 9616
rect 12310 9560 14162 9616
rect 12249 9558 14162 9560
rect 12249 9555 12315 9558
rect 13362 9528 14162 9558
rect 2922 9280 3242 9281
rect 2922 9216 2930 9280
rect 2994 9216 3010 9280
rect 3074 9216 3090 9280
rect 3154 9216 3170 9280
rect 3234 9216 3242 9280
rect 2922 9215 3242 9216
rect 6878 9280 7198 9281
rect 6878 9216 6886 9280
rect 6950 9216 6966 9280
rect 7030 9216 7046 9280
rect 7110 9216 7126 9280
rect 7190 9216 7198 9280
rect 6878 9215 7198 9216
rect 10834 9280 11154 9281
rect 10834 9216 10842 9280
rect 10906 9216 10922 9280
rect 10986 9216 11002 9280
rect 11066 9216 11082 9280
rect 11146 9216 11154 9280
rect 10834 9215 11154 9216
rect 4900 8736 5220 8737
rect 4900 8672 4908 8736
rect 4972 8672 4988 8736
rect 5052 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5220 8736
rect 4900 8671 5220 8672
rect 8856 8736 9176 8737
rect 8856 8672 8864 8736
rect 8928 8672 8944 8736
rect 9008 8672 9024 8736
rect 9088 8672 9104 8736
rect 9168 8672 9176 8736
rect 8856 8671 9176 8672
rect 2922 8192 3242 8193
rect 2922 8128 2930 8192
rect 2994 8128 3010 8192
rect 3074 8128 3090 8192
rect 3154 8128 3170 8192
rect 3234 8128 3242 8192
rect 2922 8127 3242 8128
rect 6878 8192 7198 8193
rect 6878 8128 6886 8192
rect 6950 8128 6966 8192
rect 7030 8128 7046 8192
rect 7110 8128 7126 8192
rect 7190 8128 7198 8192
rect 6878 8127 7198 8128
rect 10834 8192 11154 8193
rect 10834 8128 10842 8192
rect 10906 8128 10922 8192
rect 10986 8128 11002 8192
rect 11066 8128 11082 8192
rect 11146 8128 11154 8192
rect 10834 8127 11154 8128
rect 0 7714 800 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 800 7654
rect 1485 7651 1551 7654
rect 12249 7714 12315 7717
rect 13362 7714 14162 7744
rect 12249 7712 14162 7714
rect 12249 7656 12254 7712
rect 12310 7656 14162 7712
rect 12249 7654 14162 7656
rect 12249 7651 12315 7654
rect 4900 7648 5220 7649
rect 4900 7584 4908 7648
rect 4972 7584 4988 7648
rect 5052 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5220 7648
rect 4900 7583 5220 7584
rect 8856 7648 9176 7649
rect 8856 7584 8864 7648
rect 8928 7584 8944 7648
rect 9008 7584 9024 7648
rect 9088 7584 9104 7648
rect 9168 7584 9176 7648
rect 13362 7624 14162 7654
rect 8856 7583 9176 7584
rect 7598 7108 7604 7172
rect 7668 7170 7674 7172
rect 7741 7170 7807 7173
rect 7668 7168 7807 7170
rect 7668 7112 7746 7168
rect 7802 7112 7807 7168
rect 7668 7110 7807 7112
rect 7668 7108 7674 7110
rect 7741 7107 7807 7110
rect 2922 7104 3242 7105
rect 2922 7040 2930 7104
rect 2994 7040 3010 7104
rect 3074 7040 3090 7104
rect 3154 7040 3170 7104
rect 3234 7040 3242 7104
rect 2922 7039 3242 7040
rect 6878 7104 7198 7105
rect 6878 7040 6886 7104
rect 6950 7040 6966 7104
rect 7030 7040 7046 7104
rect 7110 7040 7126 7104
rect 7190 7040 7198 7104
rect 6878 7039 7198 7040
rect 10834 7104 11154 7105
rect 10834 7040 10842 7104
rect 10906 7040 10922 7104
rect 10986 7040 11002 7104
rect 11066 7040 11082 7104
rect 11146 7040 11154 7104
rect 10834 7039 11154 7040
rect 7097 6898 7163 6901
rect 8845 6898 8911 6901
rect 7097 6896 8911 6898
rect 7097 6840 7102 6896
rect 7158 6840 8850 6896
rect 8906 6840 8911 6896
rect 7097 6838 8911 6840
rect 7097 6835 7163 6838
rect 8845 6835 8911 6838
rect 2405 6762 2471 6765
rect 12065 6762 12131 6765
rect 2405 6760 12131 6762
rect 2405 6704 2410 6760
rect 2466 6704 12070 6760
rect 12126 6704 12131 6760
rect 2405 6702 12131 6704
rect 2405 6699 2471 6702
rect 12065 6699 12131 6702
rect 9673 6624 9739 6629
rect 9857 6626 9923 6629
rect 9673 6568 9678 6624
rect 9734 6568 9739 6624
rect 9673 6563 9739 6568
rect 9814 6624 9923 6626
rect 9814 6568 9862 6624
rect 9918 6568 9923 6624
rect 9814 6563 9923 6568
rect 4900 6560 5220 6561
rect 4900 6496 4908 6560
rect 4972 6496 4988 6560
rect 5052 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5220 6560
rect 4900 6495 5220 6496
rect 8856 6560 9176 6561
rect 8856 6496 8864 6560
rect 8928 6496 8944 6560
rect 9008 6496 9024 6560
rect 9088 6496 9104 6560
rect 9168 6496 9176 6560
rect 8856 6495 9176 6496
rect 7189 6490 7255 6493
rect 8569 6490 8635 6493
rect 7189 6488 8635 6490
rect 7189 6432 7194 6488
rect 7250 6432 8574 6488
rect 8630 6432 8635 6488
rect 7189 6430 8635 6432
rect 7189 6427 7255 6430
rect 8569 6427 8635 6430
rect 4429 6354 4495 6357
rect 6729 6354 6795 6357
rect 4429 6352 6795 6354
rect 4429 6296 4434 6352
rect 4490 6296 6734 6352
rect 6790 6296 6795 6352
rect 4429 6294 6795 6296
rect 4429 6291 4495 6294
rect 6729 6291 6795 6294
rect 4429 6218 4495 6221
rect 9029 6218 9095 6221
rect 4429 6216 9095 6218
rect 4429 6160 4434 6216
rect 4490 6160 9034 6216
rect 9090 6160 9095 6216
rect 4429 6158 9095 6160
rect 4429 6155 4495 6158
rect 9029 6155 9095 6158
rect 2922 6016 3242 6017
rect 2922 5952 2930 6016
rect 2994 5952 3010 6016
rect 3074 5952 3090 6016
rect 3154 5952 3170 6016
rect 3234 5952 3242 6016
rect 2922 5951 3242 5952
rect 6878 6016 7198 6017
rect 6878 5952 6886 6016
rect 6950 5952 6966 6016
rect 7030 5952 7046 6016
rect 7110 5952 7126 6016
rect 7190 5952 7198 6016
rect 6878 5951 7198 5952
rect 9676 5949 9736 6563
rect 9814 6221 9874 6563
rect 9949 6492 10015 6493
rect 9949 6488 9996 6492
rect 10060 6490 10066 6492
rect 9949 6432 9954 6488
rect 9949 6428 9996 6432
rect 10060 6430 10106 6490
rect 10060 6428 10066 6430
rect 9949 6427 10015 6428
rect 9949 6354 10015 6357
rect 10409 6354 10475 6357
rect 9949 6352 10475 6354
rect 9949 6296 9954 6352
rect 10010 6296 10414 6352
rect 10470 6296 10475 6352
rect 9949 6294 10475 6296
rect 9949 6291 10015 6294
rect 10409 6291 10475 6294
rect 9814 6216 9923 6221
rect 9814 6160 9862 6216
rect 9918 6160 9923 6216
rect 9814 6158 9923 6160
rect 9857 6155 9923 6158
rect 10834 6016 11154 6017
rect 10834 5952 10842 6016
rect 10906 5952 10922 6016
rect 10986 5952 11002 6016
rect 11066 5952 11082 6016
rect 11146 5952 11154 6016
rect 10834 5951 11154 5952
rect 9673 5944 9739 5949
rect 9673 5888 9678 5944
rect 9734 5888 9739 5944
rect 9673 5883 9739 5888
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 6821 5810 6887 5813
rect 10869 5810 10935 5813
rect 6821 5808 10935 5810
rect 6821 5752 6826 5808
rect 6882 5752 10874 5808
rect 10930 5752 10935 5808
rect 6821 5750 10935 5752
rect 6821 5747 6887 5750
rect 10869 5747 10935 5750
rect 12157 5810 12223 5813
rect 13362 5810 14162 5840
rect 12157 5808 14162 5810
rect 12157 5752 12162 5808
rect 12218 5752 14162 5808
rect 12157 5750 14162 5752
rect 12157 5747 12223 5750
rect 13362 5720 14162 5750
rect 7557 5676 7623 5677
rect 7557 5674 7604 5676
rect 7512 5672 7604 5674
rect 7668 5674 7674 5676
rect 11513 5674 11579 5677
rect 7668 5672 11579 5674
rect 7512 5616 7562 5672
rect 7668 5616 11518 5672
rect 11574 5616 11579 5672
rect 7512 5614 7604 5616
rect 7557 5612 7604 5614
rect 7668 5614 11579 5616
rect 7668 5612 7674 5614
rect 7557 5611 7623 5612
rect 11513 5611 11579 5614
rect 10225 5538 10291 5541
rect 10777 5538 10843 5541
rect 10225 5536 10843 5538
rect 10225 5480 10230 5536
rect 10286 5480 10782 5536
rect 10838 5480 10843 5536
rect 10225 5478 10843 5480
rect 10225 5475 10291 5478
rect 10777 5475 10843 5478
rect 4900 5472 5220 5473
rect 4900 5408 4908 5472
rect 4972 5408 4988 5472
rect 5052 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5220 5472
rect 4900 5407 5220 5408
rect 8856 5472 9176 5473
rect 8856 5408 8864 5472
rect 8928 5408 8944 5472
rect 9008 5408 9024 5472
rect 9088 5408 9104 5472
rect 9168 5408 9176 5472
rect 8856 5407 9176 5408
rect 9765 5402 9831 5405
rect 11881 5402 11947 5405
rect 9765 5400 11947 5402
rect 9765 5344 9770 5400
rect 9826 5344 11886 5400
rect 11942 5344 11947 5400
rect 9765 5342 11947 5344
rect 9765 5339 9831 5342
rect 11881 5339 11947 5342
rect 5809 5266 5875 5269
rect 9581 5266 9647 5269
rect 5809 5264 9647 5266
rect 5809 5208 5814 5264
rect 5870 5208 9586 5264
rect 9642 5208 9647 5264
rect 5809 5206 9647 5208
rect 5809 5203 5875 5206
rect 9581 5203 9647 5206
rect 10133 5266 10199 5269
rect 11973 5266 12039 5269
rect 10133 5264 12039 5266
rect 10133 5208 10138 5264
rect 10194 5208 11978 5264
rect 12034 5208 12039 5264
rect 10133 5206 12039 5208
rect 10133 5203 10199 5206
rect 11973 5203 12039 5206
rect 2922 4928 3242 4929
rect 2922 4864 2930 4928
rect 2994 4864 3010 4928
rect 3074 4864 3090 4928
rect 3154 4864 3170 4928
rect 3234 4864 3242 4928
rect 2922 4863 3242 4864
rect 6878 4928 7198 4929
rect 6878 4864 6886 4928
rect 6950 4864 6966 4928
rect 7030 4864 7046 4928
rect 7110 4864 7126 4928
rect 7190 4864 7198 4928
rect 6878 4863 7198 4864
rect 10834 4928 11154 4929
rect 10834 4864 10842 4928
rect 10906 4864 10922 4928
rect 10986 4864 11002 4928
rect 11066 4864 11082 4928
rect 11146 4864 11154 4928
rect 10834 4863 11154 4864
rect 4900 4384 5220 4385
rect 4900 4320 4908 4384
rect 4972 4320 4988 4384
rect 5052 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5220 4384
rect 4900 4319 5220 4320
rect 8856 4384 9176 4385
rect 8856 4320 8864 4384
rect 8928 4320 8944 4384
rect 9008 4320 9024 4384
rect 9088 4320 9104 4384
rect 9168 4320 9176 4384
rect 8856 4319 9176 4320
rect 9949 4044 10015 4045
rect 9949 4042 9996 4044
rect 9904 4040 9996 4042
rect 9904 3984 9954 4040
rect 9904 3982 9996 3984
rect 9949 3980 9996 3982
rect 10060 3980 10066 4044
rect 9949 3979 10015 3980
rect 0 3906 800 3936
rect 1853 3906 1919 3909
rect 0 3904 1919 3906
rect 0 3848 1858 3904
rect 1914 3848 1919 3904
rect 0 3846 1919 3848
rect 0 3816 800 3846
rect 1853 3843 1919 3846
rect 12157 3906 12223 3909
rect 13362 3906 14162 3936
rect 12157 3904 14162 3906
rect 12157 3848 12162 3904
rect 12218 3848 14162 3904
rect 12157 3846 14162 3848
rect 12157 3843 12223 3846
rect 2922 3840 3242 3841
rect 2922 3776 2930 3840
rect 2994 3776 3010 3840
rect 3074 3776 3090 3840
rect 3154 3776 3170 3840
rect 3234 3776 3242 3840
rect 2922 3775 3242 3776
rect 6878 3840 7198 3841
rect 6878 3776 6886 3840
rect 6950 3776 6966 3840
rect 7030 3776 7046 3840
rect 7110 3776 7126 3840
rect 7190 3776 7198 3840
rect 6878 3775 7198 3776
rect 10834 3840 11154 3841
rect 10834 3776 10842 3840
rect 10906 3776 10922 3840
rect 10986 3776 11002 3840
rect 11066 3776 11082 3840
rect 11146 3776 11154 3840
rect 13362 3816 14162 3846
rect 10834 3775 11154 3776
rect 4900 3296 5220 3297
rect 4900 3232 4908 3296
rect 4972 3232 4988 3296
rect 5052 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5220 3296
rect 4900 3231 5220 3232
rect 8856 3296 9176 3297
rect 8856 3232 8864 3296
rect 8928 3232 8944 3296
rect 9008 3232 9024 3296
rect 9088 3232 9104 3296
rect 9168 3232 9176 3296
rect 8856 3231 9176 3232
rect 2922 2752 3242 2753
rect 2922 2688 2930 2752
rect 2994 2688 3010 2752
rect 3074 2688 3090 2752
rect 3154 2688 3170 2752
rect 3234 2688 3242 2752
rect 2922 2687 3242 2688
rect 6878 2752 7198 2753
rect 6878 2688 6886 2752
rect 6950 2688 6966 2752
rect 7030 2688 7046 2752
rect 7110 2688 7126 2752
rect 7190 2688 7198 2752
rect 6878 2687 7198 2688
rect 10834 2752 11154 2753
rect 10834 2688 10842 2752
rect 10906 2688 10922 2752
rect 10986 2688 11002 2752
rect 11066 2688 11082 2752
rect 11146 2688 11154 2752
rect 10834 2687 11154 2688
rect 4900 2208 5220 2209
rect 4900 2144 4908 2208
rect 4972 2144 4988 2208
rect 5052 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5220 2208
rect 4900 2143 5220 2144
rect 8856 2208 9176 2209
rect 8856 2144 8864 2208
rect 8928 2144 8944 2208
rect 9008 2144 9024 2208
rect 9088 2144 9104 2208
rect 9168 2144 9176 2208
rect 8856 2143 9176 2144
rect 0 2002 800 2032
rect 1393 2002 1459 2005
rect 0 2000 1459 2002
rect 0 1944 1398 2000
rect 1454 1944 1459 2000
rect 0 1942 1459 1944
rect 0 1912 800 1942
rect 1393 1939 1459 1942
rect 10409 2002 10475 2005
rect 13362 2002 14162 2032
rect 10409 2000 14162 2002
rect 10409 1944 10414 2000
rect 10470 1944 14162 2000
rect 10409 1942 14162 1944
rect 10409 1939 10475 1942
rect 13362 1912 14162 1942
rect 9673 98 9739 101
rect 13362 98 14162 128
rect 9673 96 14162 98
rect 9673 40 9678 96
rect 9734 40 14162 96
rect 9673 38 14162 40
rect 9673 35 9739 38
rect 13362 8 14162 38
<< via3 >>
rect 2930 13628 2994 13632
rect 2930 13572 2934 13628
rect 2934 13572 2990 13628
rect 2990 13572 2994 13628
rect 2930 13568 2994 13572
rect 3010 13628 3074 13632
rect 3010 13572 3014 13628
rect 3014 13572 3070 13628
rect 3070 13572 3074 13628
rect 3010 13568 3074 13572
rect 3090 13628 3154 13632
rect 3090 13572 3094 13628
rect 3094 13572 3150 13628
rect 3150 13572 3154 13628
rect 3090 13568 3154 13572
rect 3170 13628 3234 13632
rect 3170 13572 3174 13628
rect 3174 13572 3230 13628
rect 3230 13572 3234 13628
rect 3170 13568 3234 13572
rect 6886 13628 6950 13632
rect 6886 13572 6890 13628
rect 6890 13572 6946 13628
rect 6946 13572 6950 13628
rect 6886 13568 6950 13572
rect 6966 13628 7030 13632
rect 6966 13572 6970 13628
rect 6970 13572 7026 13628
rect 7026 13572 7030 13628
rect 6966 13568 7030 13572
rect 7046 13628 7110 13632
rect 7046 13572 7050 13628
rect 7050 13572 7106 13628
rect 7106 13572 7110 13628
rect 7046 13568 7110 13572
rect 7126 13628 7190 13632
rect 7126 13572 7130 13628
rect 7130 13572 7186 13628
rect 7186 13572 7190 13628
rect 7126 13568 7190 13572
rect 10842 13628 10906 13632
rect 10842 13572 10846 13628
rect 10846 13572 10902 13628
rect 10902 13572 10906 13628
rect 10842 13568 10906 13572
rect 10922 13628 10986 13632
rect 10922 13572 10926 13628
rect 10926 13572 10982 13628
rect 10982 13572 10986 13628
rect 10922 13568 10986 13572
rect 11002 13628 11066 13632
rect 11002 13572 11006 13628
rect 11006 13572 11062 13628
rect 11062 13572 11066 13628
rect 11002 13568 11066 13572
rect 11082 13628 11146 13632
rect 11082 13572 11086 13628
rect 11086 13572 11142 13628
rect 11142 13572 11146 13628
rect 11082 13568 11146 13572
rect 4908 13084 4972 13088
rect 4908 13028 4912 13084
rect 4912 13028 4968 13084
rect 4968 13028 4972 13084
rect 4908 13024 4972 13028
rect 4988 13084 5052 13088
rect 4988 13028 4992 13084
rect 4992 13028 5048 13084
rect 5048 13028 5052 13084
rect 4988 13024 5052 13028
rect 5068 13084 5132 13088
rect 5068 13028 5072 13084
rect 5072 13028 5128 13084
rect 5128 13028 5132 13084
rect 5068 13024 5132 13028
rect 5148 13084 5212 13088
rect 5148 13028 5152 13084
rect 5152 13028 5208 13084
rect 5208 13028 5212 13084
rect 5148 13024 5212 13028
rect 8864 13084 8928 13088
rect 8864 13028 8868 13084
rect 8868 13028 8924 13084
rect 8924 13028 8928 13084
rect 8864 13024 8928 13028
rect 8944 13084 9008 13088
rect 8944 13028 8948 13084
rect 8948 13028 9004 13084
rect 9004 13028 9008 13084
rect 8944 13024 9008 13028
rect 9024 13084 9088 13088
rect 9024 13028 9028 13084
rect 9028 13028 9084 13084
rect 9084 13028 9088 13084
rect 9024 13024 9088 13028
rect 9104 13084 9168 13088
rect 9104 13028 9108 13084
rect 9108 13028 9164 13084
rect 9164 13028 9168 13084
rect 9104 13024 9168 13028
rect 2930 12540 2994 12544
rect 2930 12484 2934 12540
rect 2934 12484 2990 12540
rect 2990 12484 2994 12540
rect 2930 12480 2994 12484
rect 3010 12540 3074 12544
rect 3010 12484 3014 12540
rect 3014 12484 3070 12540
rect 3070 12484 3074 12540
rect 3010 12480 3074 12484
rect 3090 12540 3154 12544
rect 3090 12484 3094 12540
rect 3094 12484 3150 12540
rect 3150 12484 3154 12540
rect 3090 12480 3154 12484
rect 3170 12540 3234 12544
rect 3170 12484 3174 12540
rect 3174 12484 3230 12540
rect 3230 12484 3234 12540
rect 3170 12480 3234 12484
rect 6886 12540 6950 12544
rect 6886 12484 6890 12540
rect 6890 12484 6946 12540
rect 6946 12484 6950 12540
rect 6886 12480 6950 12484
rect 6966 12540 7030 12544
rect 6966 12484 6970 12540
rect 6970 12484 7026 12540
rect 7026 12484 7030 12540
rect 6966 12480 7030 12484
rect 7046 12540 7110 12544
rect 7046 12484 7050 12540
rect 7050 12484 7106 12540
rect 7106 12484 7110 12540
rect 7046 12480 7110 12484
rect 7126 12540 7190 12544
rect 7126 12484 7130 12540
rect 7130 12484 7186 12540
rect 7186 12484 7190 12540
rect 7126 12480 7190 12484
rect 10842 12540 10906 12544
rect 10842 12484 10846 12540
rect 10846 12484 10902 12540
rect 10902 12484 10906 12540
rect 10842 12480 10906 12484
rect 10922 12540 10986 12544
rect 10922 12484 10926 12540
rect 10926 12484 10982 12540
rect 10982 12484 10986 12540
rect 10922 12480 10986 12484
rect 11002 12540 11066 12544
rect 11002 12484 11006 12540
rect 11006 12484 11062 12540
rect 11062 12484 11066 12540
rect 11002 12480 11066 12484
rect 11082 12540 11146 12544
rect 11082 12484 11086 12540
rect 11086 12484 11142 12540
rect 11142 12484 11146 12540
rect 11082 12480 11146 12484
rect 4908 11996 4972 12000
rect 4908 11940 4912 11996
rect 4912 11940 4968 11996
rect 4968 11940 4972 11996
rect 4908 11936 4972 11940
rect 4988 11996 5052 12000
rect 4988 11940 4992 11996
rect 4992 11940 5048 11996
rect 5048 11940 5052 11996
rect 4988 11936 5052 11940
rect 5068 11996 5132 12000
rect 5068 11940 5072 11996
rect 5072 11940 5128 11996
rect 5128 11940 5132 11996
rect 5068 11936 5132 11940
rect 5148 11996 5212 12000
rect 5148 11940 5152 11996
rect 5152 11940 5208 11996
rect 5208 11940 5212 11996
rect 5148 11936 5212 11940
rect 8864 11996 8928 12000
rect 8864 11940 8868 11996
rect 8868 11940 8924 11996
rect 8924 11940 8928 11996
rect 8864 11936 8928 11940
rect 8944 11996 9008 12000
rect 8944 11940 8948 11996
rect 8948 11940 9004 11996
rect 9004 11940 9008 11996
rect 8944 11936 9008 11940
rect 9024 11996 9088 12000
rect 9024 11940 9028 11996
rect 9028 11940 9084 11996
rect 9084 11940 9088 11996
rect 9024 11936 9088 11940
rect 9104 11996 9168 12000
rect 9104 11940 9108 11996
rect 9108 11940 9164 11996
rect 9164 11940 9168 11996
rect 9104 11936 9168 11940
rect 2930 11452 2994 11456
rect 2930 11396 2934 11452
rect 2934 11396 2990 11452
rect 2990 11396 2994 11452
rect 2930 11392 2994 11396
rect 3010 11452 3074 11456
rect 3010 11396 3014 11452
rect 3014 11396 3070 11452
rect 3070 11396 3074 11452
rect 3010 11392 3074 11396
rect 3090 11452 3154 11456
rect 3090 11396 3094 11452
rect 3094 11396 3150 11452
rect 3150 11396 3154 11452
rect 3090 11392 3154 11396
rect 3170 11452 3234 11456
rect 3170 11396 3174 11452
rect 3174 11396 3230 11452
rect 3230 11396 3234 11452
rect 3170 11392 3234 11396
rect 6886 11452 6950 11456
rect 6886 11396 6890 11452
rect 6890 11396 6946 11452
rect 6946 11396 6950 11452
rect 6886 11392 6950 11396
rect 6966 11452 7030 11456
rect 6966 11396 6970 11452
rect 6970 11396 7026 11452
rect 7026 11396 7030 11452
rect 6966 11392 7030 11396
rect 7046 11452 7110 11456
rect 7046 11396 7050 11452
rect 7050 11396 7106 11452
rect 7106 11396 7110 11452
rect 7046 11392 7110 11396
rect 7126 11452 7190 11456
rect 7126 11396 7130 11452
rect 7130 11396 7186 11452
rect 7186 11396 7190 11452
rect 7126 11392 7190 11396
rect 10842 11452 10906 11456
rect 10842 11396 10846 11452
rect 10846 11396 10902 11452
rect 10902 11396 10906 11452
rect 10842 11392 10906 11396
rect 10922 11452 10986 11456
rect 10922 11396 10926 11452
rect 10926 11396 10982 11452
rect 10982 11396 10986 11452
rect 10922 11392 10986 11396
rect 11002 11452 11066 11456
rect 11002 11396 11006 11452
rect 11006 11396 11062 11452
rect 11062 11396 11066 11452
rect 11002 11392 11066 11396
rect 11082 11452 11146 11456
rect 11082 11396 11086 11452
rect 11086 11396 11142 11452
rect 11142 11396 11146 11452
rect 11082 11392 11146 11396
rect 4908 10908 4972 10912
rect 4908 10852 4912 10908
rect 4912 10852 4968 10908
rect 4968 10852 4972 10908
rect 4908 10848 4972 10852
rect 4988 10908 5052 10912
rect 4988 10852 4992 10908
rect 4992 10852 5048 10908
rect 5048 10852 5052 10908
rect 4988 10848 5052 10852
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 8864 10908 8928 10912
rect 8864 10852 8868 10908
rect 8868 10852 8924 10908
rect 8924 10852 8928 10908
rect 8864 10848 8928 10852
rect 8944 10908 9008 10912
rect 8944 10852 8948 10908
rect 8948 10852 9004 10908
rect 9004 10852 9008 10908
rect 8944 10848 9008 10852
rect 9024 10908 9088 10912
rect 9024 10852 9028 10908
rect 9028 10852 9084 10908
rect 9084 10852 9088 10908
rect 9024 10848 9088 10852
rect 9104 10908 9168 10912
rect 9104 10852 9108 10908
rect 9108 10852 9164 10908
rect 9164 10852 9168 10908
rect 9104 10848 9168 10852
rect 2930 10364 2994 10368
rect 2930 10308 2934 10364
rect 2934 10308 2990 10364
rect 2990 10308 2994 10364
rect 2930 10304 2994 10308
rect 3010 10364 3074 10368
rect 3010 10308 3014 10364
rect 3014 10308 3070 10364
rect 3070 10308 3074 10364
rect 3010 10304 3074 10308
rect 3090 10364 3154 10368
rect 3090 10308 3094 10364
rect 3094 10308 3150 10364
rect 3150 10308 3154 10364
rect 3090 10304 3154 10308
rect 3170 10364 3234 10368
rect 3170 10308 3174 10364
rect 3174 10308 3230 10364
rect 3230 10308 3234 10364
rect 3170 10304 3234 10308
rect 6886 10364 6950 10368
rect 6886 10308 6890 10364
rect 6890 10308 6946 10364
rect 6946 10308 6950 10364
rect 6886 10304 6950 10308
rect 6966 10364 7030 10368
rect 6966 10308 6970 10364
rect 6970 10308 7026 10364
rect 7026 10308 7030 10364
rect 6966 10304 7030 10308
rect 7046 10364 7110 10368
rect 7046 10308 7050 10364
rect 7050 10308 7106 10364
rect 7106 10308 7110 10364
rect 7046 10304 7110 10308
rect 7126 10364 7190 10368
rect 7126 10308 7130 10364
rect 7130 10308 7186 10364
rect 7186 10308 7190 10364
rect 7126 10304 7190 10308
rect 10842 10364 10906 10368
rect 10842 10308 10846 10364
rect 10846 10308 10902 10364
rect 10902 10308 10906 10364
rect 10842 10304 10906 10308
rect 10922 10364 10986 10368
rect 10922 10308 10926 10364
rect 10926 10308 10982 10364
rect 10982 10308 10986 10364
rect 10922 10304 10986 10308
rect 11002 10364 11066 10368
rect 11002 10308 11006 10364
rect 11006 10308 11062 10364
rect 11062 10308 11066 10364
rect 11002 10304 11066 10308
rect 11082 10364 11146 10368
rect 11082 10308 11086 10364
rect 11086 10308 11142 10364
rect 11142 10308 11146 10364
rect 11082 10304 11146 10308
rect 4908 9820 4972 9824
rect 4908 9764 4912 9820
rect 4912 9764 4968 9820
rect 4968 9764 4972 9820
rect 4908 9760 4972 9764
rect 4988 9820 5052 9824
rect 4988 9764 4992 9820
rect 4992 9764 5048 9820
rect 5048 9764 5052 9820
rect 4988 9760 5052 9764
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 8864 9820 8928 9824
rect 8864 9764 8868 9820
rect 8868 9764 8924 9820
rect 8924 9764 8928 9820
rect 8864 9760 8928 9764
rect 8944 9820 9008 9824
rect 8944 9764 8948 9820
rect 8948 9764 9004 9820
rect 9004 9764 9008 9820
rect 8944 9760 9008 9764
rect 9024 9820 9088 9824
rect 9024 9764 9028 9820
rect 9028 9764 9084 9820
rect 9084 9764 9088 9820
rect 9024 9760 9088 9764
rect 9104 9820 9168 9824
rect 9104 9764 9108 9820
rect 9108 9764 9164 9820
rect 9164 9764 9168 9820
rect 9104 9760 9168 9764
rect 2930 9276 2994 9280
rect 2930 9220 2934 9276
rect 2934 9220 2990 9276
rect 2990 9220 2994 9276
rect 2930 9216 2994 9220
rect 3010 9276 3074 9280
rect 3010 9220 3014 9276
rect 3014 9220 3070 9276
rect 3070 9220 3074 9276
rect 3010 9216 3074 9220
rect 3090 9276 3154 9280
rect 3090 9220 3094 9276
rect 3094 9220 3150 9276
rect 3150 9220 3154 9276
rect 3090 9216 3154 9220
rect 3170 9276 3234 9280
rect 3170 9220 3174 9276
rect 3174 9220 3230 9276
rect 3230 9220 3234 9276
rect 3170 9216 3234 9220
rect 6886 9276 6950 9280
rect 6886 9220 6890 9276
rect 6890 9220 6946 9276
rect 6946 9220 6950 9276
rect 6886 9216 6950 9220
rect 6966 9276 7030 9280
rect 6966 9220 6970 9276
rect 6970 9220 7026 9276
rect 7026 9220 7030 9276
rect 6966 9216 7030 9220
rect 7046 9276 7110 9280
rect 7046 9220 7050 9276
rect 7050 9220 7106 9276
rect 7106 9220 7110 9276
rect 7046 9216 7110 9220
rect 7126 9276 7190 9280
rect 7126 9220 7130 9276
rect 7130 9220 7186 9276
rect 7186 9220 7190 9276
rect 7126 9216 7190 9220
rect 10842 9276 10906 9280
rect 10842 9220 10846 9276
rect 10846 9220 10902 9276
rect 10902 9220 10906 9276
rect 10842 9216 10906 9220
rect 10922 9276 10986 9280
rect 10922 9220 10926 9276
rect 10926 9220 10982 9276
rect 10982 9220 10986 9276
rect 10922 9216 10986 9220
rect 11002 9276 11066 9280
rect 11002 9220 11006 9276
rect 11006 9220 11062 9276
rect 11062 9220 11066 9276
rect 11002 9216 11066 9220
rect 11082 9276 11146 9280
rect 11082 9220 11086 9276
rect 11086 9220 11142 9276
rect 11142 9220 11146 9276
rect 11082 9216 11146 9220
rect 4908 8732 4972 8736
rect 4908 8676 4912 8732
rect 4912 8676 4968 8732
rect 4968 8676 4972 8732
rect 4908 8672 4972 8676
rect 4988 8732 5052 8736
rect 4988 8676 4992 8732
rect 4992 8676 5048 8732
rect 5048 8676 5052 8732
rect 4988 8672 5052 8676
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 8864 8732 8928 8736
rect 8864 8676 8868 8732
rect 8868 8676 8924 8732
rect 8924 8676 8928 8732
rect 8864 8672 8928 8676
rect 8944 8732 9008 8736
rect 8944 8676 8948 8732
rect 8948 8676 9004 8732
rect 9004 8676 9008 8732
rect 8944 8672 9008 8676
rect 9024 8732 9088 8736
rect 9024 8676 9028 8732
rect 9028 8676 9084 8732
rect 9084 8676 9088 8732
rect 9024 8672 9088 8676
rect 9104 8732 9168 8736
rect 9104 8676 9108 8732
rect 9108 8676 9164 8732
rect 9164 8676 9168 8732
rect 9104 8672 9168 8676
rect 2930 8188 2994 8192
rect 2930 8132 2934 8188
rect 2934 8132 2990 8188
rect 2990 8132 2994 8188
rect 2930 8128 2994 8132
rect 3010 8188 3074 8192
rect 3010 8132 3014 8188
rect 3014 8132 3070 8188
rect 3070 8132 3074 8188
rect 3010 8128 3074 8132
rect 3090 8188 3154 8192
rect 3090 8132 3094 8188
rect 3094 8132 3150 8188
rect 3150 8132 3154 8188
rect 3090 8128 3154 8132
rect 3170 8188 3234 8192
rect 3170 8132 3174 8188
rect 3174 8132 3230 8188
rect 3230 8132 3234 8188
rect 3170 8128 3234 8132
rect 6886 8188 6950 8192
rect 6886 8132 6890 8188
rect 6890 8132 6946 8188
rect 6946 8132 6950 8188
rect 6886 8128 6950 8132
rect 6966 8188 7030 8192
rect 6966 8132 6970 8188
rect 6970 8132 7026 8188
rect 7026 8132 7030 8188
rect 6966 8128 7030 8132
rect 7046 8188 7110 8192
rect 7046 8132 7050 8188
rect 7050 8132 7106 8188
rect 7106 8132 7110 8188
rect 7046 8128 7110 8132
rect 7126 8188 7190 8192
rect 7126 8132 7130 8188
rect 7130 8132 7186 8188
rect 7186 8132 7190 8188
rect 7126 8128 7190 8132
rect 10842 8188 10906 8192
rect 10842 8132 10846 8188
rect 10846 8132 10902 8188
rect 10902 8132 10906 8188
rect 10842 8128 10906 8132
rect 10922 8188 10986 8192
rect 10922 8132 10926 8188
rect 10926 8132 10982 8188
rect 10982 8132 10986 8188
rect 10922 8128 10986 8132
rect 11002 8188 11066 8192
rect 11002 8132 11006 8188
rect 11006 8132 11062 8188
rect 11062 8132 11066 8188
rect 11002 8128 11066 8132
rect 11082 8188 11146 8192
rect 11082 8132 11086 8188
rect 11086 8132 11142 8188
rect 11142 8132 11146 8188
rect 11082 8128 11146 8132
rect 4908 7644 4972 7648
rect 4908 7588 4912 7644
rect 4912 7588 4968 7644
rect 4968 7588 4972 7644
rect 4908 7584 4972 7588
rect 4988 7644 5052 7648
rect 4988 7588 4992 7644
rect 4992 7588 5048 7644
rect 5048 7588 5052 7644
rect 4988 7584 5052 7588
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 8864 7644 8928 7648
rect 8864 7588 8868 7644
rect 8868 7588 8924 7644
rect 8924 7588 8928 7644
rect 8864 7584 8928 7588
rect 8944 7644 9008 7648
rect 8944 7588 8948 7644
rect 8948 7588 9004 7644
rect 9004 7588 9008 7644
rect 8944 7584 9008 7588
rect 9024 7644 9088 7648
rect 9024 7588 9028 7644
rect 9028 7588 9084 7644
rect 9084 7588 9088 7644
rect 9024 7584 9088 7588
rect 9104 7644 9168 7648
rect 9104 7588 9108 7644
rect 9108 7588 9164 7644
rect 9164 7588 9168 7644
rect 9104 7584 9168 7588
rect 7604 7108 7668 7172
rect 2930 7100 2994 7104
rect 2930 7044 2934 7100
rect 2934 7044 2990 7100
rect 2990 7044 2994 7100
rect 2930 7040 2994 7044
rect 3010 7100 3074 7104
rect 3010 7044 3014 7100
rect 3014 7044 3070 7100
rect 3070 7044 3074 7100
rect 3010 7040 3074 7044
rect 3090 7100 3154 7104
rect 3090 7044 3094 7100
rect 3094 7044 3150 7100
rect 3150 7044 3154 7100
rect 3090 7040 3154 7044
rect 3170 7100 3234 7104
rect 3170 7044 3174 7100
rect 3174 7044 3230 7100
rect 3230 7044 3234 7100
rect 3170 7040 3234 7044
rect 6886 7100 6950 7104
rect 6886 7044 6890 7100
rect 6890 7044 6946 7100
rect 6946 7044 6950 7100
rect 6886 7040 6950 7044
rect 6966 7100 7030 7104
rect 6966 7044 6970 7100
rect 6970 7044 7026 7100
rect 7026 7044 7030 7100
rect 6966 7040 7030 7044
rect 7046 7100 7110 7104
rect 7046 7044 7050 7100
rect 7050 7044 7106 7100
rect 7106 7044 7110 7100
rect 7046 7040 7110 7044
rect 7126 7100 7190 7104
rect 7126 7044 7130 7100
rect 7130 7044 7186 7100
rect 7186 7044 7190 7100
rect 7126 7040 7190 7044
rect 10842 7100 10906 7104
rect 10842 7044 10846 7100
rect 10846 7044 10902 7100
rect 10902 7044 10906 7100
rect 10842 7040 10906 7044
rect 10922 7100 10986 7104
rect 10922 7044 10926 7100
rect 10926 7044 10982 7100
rect 10982 7044 10986 7100
rect 10922 7040 10986 7044
rect 11002 7100 11066 7104
rect 11002 7044 11006 7100
rect 11006 7044 11062 7100
rect 11062 7044 11066 7100
rect 11002 7040 11066 7044
rect 11082 7100 11146 7104
rect 11082 7044 11086 7100
rect 11086 7044 11142 7100
rect 11142 7044 11146 7100
rect 11082 7040 11146 7044
rect 4908 6556 4972 6560
rect 4908 6500 4912 6556
rect 4912 6500 4968 6556
rect 4968 6500 4972 6556
rect 4908 6496 4972 6500
rect 4988 6556 5052 6560
rect 4988 6500 4992 6556
rect 4992 6500 5048 6556
rect 5048 6500 5052 6556
rect 4988 6496 5052 6500
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 8864 6556 8928 6560
rect 8864 6500 8868 6556
rect 8868 6500 8924 6556
rect 8924 6500 8928 6556
rect 8864 6496 8928 6500
rect 8944 6556 9008 6560
rect 8944 6500 8948 6556
rect 8948 6500 9004 6556
rect 9004 6500 9008 6556
rect 8944 6496 9008 6500
rect 9024 6556 9088 6560
rect 9024 6500 9028 6556
rect 9028 6500 9084 6556
rect 9084 6500 9088 6556
rect 9024 6496 9088 6500
rect 9104 6556 9168 6560
rect 9104 6500 9108 6556
rect 9108 6500 9164 6556
rect 9164 6500 9168 6556
rect 9104 6496 9168 6500
rect 2930 6012 2994 6016
rect 2930 5956 2934 6012
rect 2934 5956 2990 6012
rect 2990 5956 2994 6012
rect 2930 5952 2994 5956
rect 3010 6012 3074 6016
rect 3010 5956 3014 6012
rect 3014 5956 3070 6012
rect 3070 5956 3074 6012
rect 3010 5952 3074 5956
rect 3090 6012 3154 6016
rect 3090 5956 3094 6012
rect 3094 5956 3150 6012
rect 3150 5956 3154 6012
rect 3090 5952 3154 5956
rect 3170 6012 3234 6016
rect 3170 5956 3174 6012
rect 3174 5956 3230 6012
rect 3230 5956 3234 6012
rect 3170 5952 3234 5956
rect 6886 6012 6950 6016
rect 6886 5956 6890 6012
rect 6890 5956 6946 6012
rect 6946 5956 6950 6012
rect 6886 5952 6950 5956
rect 6966 6012 7030 6016
rect 6966 5956 6970 6012
rect 6970 5956 7026 6012
rect 7026 5956 7030 6012
rect 6966 5952 7030 5956
rect 7046 6012 7110 6016
rect 7046 5956 7050 6012
rect 7050 5956 7106 6012
rect 7106 5956 7110 6012
rect 7046 5952 7110 5956
rect 7126 6012 7190 6016
rect 7126 5956 7130 6012
rect 7130 5956 7186 6012
rect 7186 5956 7190 6012
rect 7126 5952 7190 5956
rect 9996 6488 10060 6492
rect 9996 6432 10010 6488
rect 10010 6432 10060 6488
rect 9996 6428 10060 6432
rect 10842 6012 10906 6016
rect 10842 5956 10846 6012
rect 10846 5956 10902 6012
rect 10902 5956 10906 6012
rect 10842 5952 10906 5956
rect 10922 6012 10986 6016
rect 10922 5956 10926 6012
rect 10926 5956 10982 6012
rect 10982 5956 10986 6012
rect 10922 5952 10986 5956
rect 11002 6012 11066 6016
rect 11002 5956 11006 6012
rect 11006 5956 11062 6012
rect 11062 5956 11066 6012
rect 11002 5952 11066 5956
rect 11082 6012 11146 6016
rect 11082 5956 11086 6012
rect 11086 5956 11142 6012
rect 11142 5956 11146 6012
rect 11082 5952 11146 5956
rect 7604 5672 7668 5676
rect 7604 5616 7618 5672
rect 7618 5616 7668 5672
rect 7604 5612 7668 5616
rect 4908 5468 4972 5472
rect 4908 5412 4912 5468
rect 4912 5412 4968 5468
rect 4968 5412 4972 5468
rect 4908 5408 4972 5412
rect 4988 5468 5052 5472
rect 4988 5412 4992 5468
rect 4992 5412 5048 5468
rect 5048 5412 5052 5468
rect 4988 5408 5052 5412
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 8864 5468 8928 5472
rect 8864 5412 8868 5468
rect 8868 5412 8924 5468
rect 8924 5412 8928 5468
rect 8864 5408 8928 5412
rect 8944 5468 9008 5472
rect 8944 5412 8948 5468
rect 8948 5412 9004 5468
rect 9004 5412 9008 5468
rect 8944 5408 9008 5412
rect 9024 5468 9088 5472
rect 9024 5412 9028 5468
rect 9028 5412 9084 5468
rect 9084 5412 9088 5468
rect 9024 5408 9088 5412
rect 9104 5468 9168 5472
rect 9104 5412 9108 5468
rect 9108 5412 9164 5468
rect 9164 5412 9168 5468
rect 9104 5408 9168 5412
rect 2930 4924 2994 4928
rect 2930 4868 2934 4924
rect 2934 4868 2990 4924
rect 2990 4868 2994 4924
rect 2930 4864 2994 4868
rect 3010 4924 3074 4928
rect 3010 4868 3014 4924
rect 3014 4868 3070 4924
rect 3070 4868 3074 4924
rect 3010 4864 3074 4868
rect 3090 4924 3154 4928
rect 3090 4868 3094 4924
rect 3094 4868 3150 4924
rect 3150 4868 3154 4924
rect 3090 4864 3154 4868
rect 3170 4924 3234 4928
rect 3170 4868 3174 4924
rect 3174 4868 3230 4924
rect 3230 4868 3234 4924
rect 3170 4864 3234 4868
rect 6886 4924 6950 4928
rect 6886 4868 6890 4924
rect 6890 4868 6946 4924
rect 6946 4868 6950 4924
rect 6886 4864 6950 4868
rect 6966 4924 7030 4928
rect 6966 4868 6970 4924
rect 6970 4868 7026 4924
rect 7026 4868 7030 4924
rect 6966 4864 7030 4868
rect 7046 4924 7110 4928
rect 7046 4868 7050 4924
rect 7050 4868 7106 4924
rect 7106 4868 7110 4924
rect 7046 4864 7110 4868
rect 7126 4924 7190 4928
rect 7126 4868 7130 4924
rect 7130 4868 7186 4924
rect 7186 4868 7190 4924
rect 7126 4864 7190 4868
rect 10842 4924 10906 4928
rect 10842 4868 10846 4924
rect 10846 4868 10902 4924
rect 10902 4868 10906 4924
rect 10842 4864 10906 4868
rect 10922 4924 10986 4928
rect 10922 4868 10926 4924
rect 10926 4868 10982 4924
rect 10982 4868 10986 4924
rect 10922 4864 10986 4868
rect 11002 4924 11066 4928
rect 11002 4868 11006 4924
rect 11006 4868 11062 4924
rect 11062 4868 11066 4924
rect 11002 4864 11066 4868
rect 11082 4924 11146 4928
rect 11082 4868 11086 4924
rect 11086 4868 11142 4924
rect 11142 4868 11146 4924
rect 11082 4864 11146 4868
rect 4908 4380 4972 4384
rect 4908 4324 4912 4380
rect 4912 4324 4968 4380
rect 4968 4324 4972 4380
rect 4908 4320 4972 4324
rect 4988 4380 5052 4384
rect 4988 4324 4992 4380
rect 4992 4324 5048 4380
rect 5048 4324 5052 4380
rect 4988 4320 5052 4324
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 8864 4380 8928 4384
rect 8864 4324 8868 4380
rect 8868 4324 8924 4380
rect 8924 4324 8928 4380
rect 8864 4320 8928 4324
rect 8944 4380 9008 4384
rect 8944 4324 8948 4380
rect 8948 4324 9004 4380
rect 9004 4324 9008 4380
rect 8944 4320 9008 4324
rect 9024 4380 9088 4384
rect 9024 4324 9028 4380
rect 9028 4324 9084 4380
rect 9084 4324 9088 4380
rect 9024 4320 9088 4324
rect 9104 4380 9168 4384
rect 9104 4324 9108 4380
rect 9108 4324 9164 4380
rect 9164 4324 9168 4380
rect 9104 4320 9168 4324
rect 9996 4040 10060 4044
rect 9996 3984 10010 4040
rect 10010 3984 10060 4040
rect 9996 3980 10060 3984
rect 2930 3836 2994 3840
rect 2930 3780 2934 3836
rect 2934 3780 2990 3836
rect 2990 3780 2994 3836
rect 2930 3776 2994 3780
rect 3010 3836 3074 3840
rect 3010 3780 3014 3836
rect 3014 3780 3070 3836
rect 3070 3780 3074 3836
rect 3010 3776 3074 3780
rect 3090 3836 3154 3840
rect 3090 3780 3094 3836
rect 3094 3780 3150 3836
rect 3150 3780 3154 3836
rect 3090 3776 3154 3780
rect 3170 3836 3234 3840
rect 3170 3780 3174 3836
rect 3174 3780 3230 3836
rect 3230 3780 3234 3836
rect 3170 3776 3234 3780
rect 6886 3836 6950 3840
rect 6886 3780 6890 3836
rect 6890 3780 6946 3836
rect 6946 3780 6950 3836
rect 6886 3776 6950 3780
rect 6966 3836 7030 3840
rect 6966 3780 6970 3836
rect 6970 3780 7026 3836
rect 7026 3780 7030 3836
rect 6966 3776 7030 3780
rect 7046 3836 7110 3840
rect 7046 3780 7050 3836
rect 7050 3780 7106 3836
rect 7106 3780 7110 3836
rect 7046 3776 7110 3780
rect 7126 3836 7190 3840
rect 7126 3780 7130 3836
rect 7130 3780 7186 3836
rect 7186 3780 7190 3836
rect 7126 3776 7190 3780
rect 10842 3836 10906 3840
rect 10842 3780 10846 3836
rect 10846 3780 10902 3836
rect 10902 3780 10906 3836
rect 10842 3776 10906 3780
rect 10922 3836 10986 3840
rect 10922 3780 10926 3836
rect 10926 3780 10982 3836
rect 10982 3780 10986 3836
rect 10922 3776 10986 3780
rect 11002 3836 11066 3840
rect 11002 3780 11006 3836
rect 11006 3780 11062 3836
rect 11062 3780 11066 3836
rect 11002 3776 11066 3780
rect 11082 3836 11146 3840
rect 11082 3780 11086 3836
rect 11086 3780 11142 3836
rect 11142 3780 11146 3836
rect 11082 3776 11146 3780
rect 4908 3292 4972 3296
rect 4908 3236 4912 3292
rect 4912 3236 4968 3292
rect 4968 3236 4972 3292
rect 4908 3232 4972 3236
rect 4988 3292 5052 3296
rect 4988 3236 4992 3292
rect 4992 3236 5048 3292
rect 5048 3236 5052 3292
rect 4988 3232 5052 3236
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 8864 3292 8928 3296
rect 8864 3236 8868 3292
rect 8868 3236 8924 3292
rect 8924 3236 8928 3292
rect 8864 3232 8928 3236
rect 8944 3292 9008 3296
rect 8944 3236 8948 3292
rect 8948 3236 9004 3292
rect 9004 3236 9008 3292
rect 8944 3232 9008 3236
rect 9024 3292 9088 3296
rect 9024 3236 9028 3292
rect 9028 3236 9084 3292
rect 9084 3236 9088 3292
rect 9024 3232 9088 3236
rect 9104 3292 9168 3296
rect 9104 3236 9108 3292
rect 9108 3236 9164 3292
rect 9164 3236 9168 3292
rect 9104 3232 9168 3236
rect 2930 2748 2994 2752
rect 2930 2692 2934 2748
rect 2934 2692 2990 2748
rect 2990 2692 2994 2748
rect 2930 2688 2994 2692
rect 3010 2748 3074 2752
rect 3010 2692 3014 2748
rect 3014 2692 3070 2748
rect 3070 2692 3074 2748
rect 3010 2688 3074 2692
rect 3090 2748 3154 2752
rect 3090 2692 3094 2748
rect 3094 2692 3150 2748
rect 3150 2692 3154 2748
rect 3090 2688 3154 2692
rect 3170 2748 3234 2752
rect 3170 2692 3174 2748
rect 3174 2692 3230 2748
rect 3230 2692 3234 2748
rect 3170 2688 3234 2692
rect 6886 2748 6950 2752
rect 6886 2692 6890 2748
rect 6890 2692 6946 2748
rect 6946 2692 6950 2748
rect 6886 2688 6950 2692
rect 6966 2748 7030 2752
rect 6966 2692 6970 2748
rect 6970 2692 7026 2748
rect 7026 2692 7030 2748
rect 6966 2688 7030 2692
rect 7046 2748 7110 2752
rect 7046 2692 7050 2748
rect 7050 2692 7106 2748
rect 7106 2692 7110 2748
rect 7046 2688 7110 2692
rect 7126 2748 7190 2752
rect 7126 2692 7130 2748
rect 7130 2692 7186 2748
rect 7186 2692 7190 2748
rect 7126 2688 7190 2692
rect 10842 2748 10906 2752
rect 10842 2692 10846 2748
rect 10846 2692 10902 2748
rect 10902 2692 10906 2748
rect 10842 2688 10906 2692
rect 10922 2748 10986 2752
rect 10922 2692 10926 2748
rect 10926 2692 10982 2748
rect 10982 2692 10986 2748
rect 10922 2688 10986 2692
rect 11002 2748 11066 2752
rect 11002 2692 11006 2748
rect 11006 2692 11062 2748
rect 11062 2692 11066 2748
rect 11002 2688 11066 2692
rect 11082 2748 11146 2752
rect 11082 2692 11086 2748
rect 11086 2692 11142 2748
rect 11142 2692 11146 2748
rect 11082 2688 11146 2692
rect 4908 2204 4972 2208
rect 4908 2148 4912 2204
rect 4912 2148 4968 2204
rect 4968 2148 4972 2204
rect 4908 2144 4972 2148
rect 4988 2204 5052 2208
rect 4988 2148 4992 2204
rect 4992 2148 5048 2204
rect 5048 2148 5052 2204
rect 4988 2144 5052 2148
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 8864 2204 8928 2208
rect 8864 2148 8868 2204
rect 8868 2148 8924 2204
rect 8924 2148 8928 2204
rect 8864 2144 8928 2148
rect 8944 2204 9008 2208
rect 8944 2148 8948 2204
rect 8948 2148 9004 2204
rect 9004 2148 9008 2204
rect 8944 2144 9008 2148
rect 9024 2204 9088 2208
rect 9024 2148 9028 2204
rect 9028 2148 9084 2204
rect 9084 2148 9088 2204
rect 9024 2144 9088 2148
rect 9104 2204 9168 2208
rect 9104 2148 9108 2204
rect 9108 2148 9164 2204
rect 9164 2148 9168 2204
rect 9104 2144 9168 2148
<< metal4 >>
rect 2922 13632 3242 13648
rect 2922 13568 2930 13632
rect 2994 13568 3010 13632
rect 3074 13568 3090 13632
rect 3154 13568 3170 13632
rect 3234 13568 3242 13632
rect 2922 12544 3242 13568
rect 2922 12480 2930 12544
rect 2994 12480 3010 12544
rect 3074 12480 3090 12544
rect 3154 12480 3170 12544
rect 3234 12480 3242 12544
rect 2922 11766 3242 12480
rect 2922 11530 2964 11766
rect 3200 11530 3242 11766
rect 2922 11456 3242 11530
rect 2922 11392 2930 11456
rect 2994 11392 3010 11456
rect 3074 11392 3090 11456
rect 3154 11392 3170 11456
rect 3234 11392 3242 11456
rect 2922 10368 3242 11392
rect 2922 10304 2930 10368
rect 2994 10304 3010 10368
rect 3074 10304 3090 10368
rect 3154 10304 3170 10368
rect 3234 10304 3242 10368
rect 2922 9280 3242 10304
rect 2922 9216 2930 9280
rect 2994 9216 3010 9280
rect 3074 9216 3090 9280
rect 3154 9216 3170 9280
rect 3234 9216 3242 9280
rect 2922 8192 3242 9216
rect 2922 8128 2930 8192
rect 2994 8128 3010 8192
rect 3074 8128 3090 8192
rect 3154 8128 3170 8192
rect 3234 8128 3242 8192
rect 2922 7958 3242 8128
rect 2922 7722 2964 7958
rect 3200 7722 3242 7958
rect 2922 7104 3242 7722
rect 2922 7040 2930 7104
rect 2994 7040 3010 7104
rect 3074 7040 3090 7104
rect 3154 7040 3170 7104
rect 3234 7040 3242 7104
rect 2922 6016 3242 7040
rect 2922 5952 2930 6016
rect 2994 5952 3010 6016
rect 3074 5952 3090 6016
rect 3154 5952 3170 6016
rect 3234 5952 3242 6016
rect 2922 4928 3242 5952
rect 2922 4864 2930 4928
rect 2994 4864 3010 4928
rect 3074 4864 3090 4928
rect 3154 4864 3170 4928
rect 3234 4864 3242 4928
rect 2922 4150 3242 4864
rect 2922 3914 2964 4150
rect 3200 3914 3242 4150
rect 2922 3840 3242 3914
rect 2922 3776 2930 3840
rect 2994 3776 3010 3840
rect 3074 3776 3090 3840
rect 3154 3776 3170 3840
rect 3234 3776 3242 3840
rect 2922 2752 3242 3776
rect 2922 2688 2930 2752
rect 2994 2688 3010 2752
rect 3074 2688 3090 2752
rect 3154 2688 3170 2752
rect 3234 2688 3242 2752
rect 2922 2128 3242 2688
rect 4900 13088 5220 13648
rect 4900 13024 4908 13088
rect 4972 13024 4988 13088
rect 5052 13024 5068 13088
rect 5132 13024 5148 13088
rect 5212 13024 5220 13088
rect 4900 12000 5220 13024
rect 4900 11936 4908 12000
rect 4972 11936 4988 12000
rect 5052 11936 5068 12000
rect 5132 11936 5148 12000
rect 5212 11936 5220 12000
rect 4900 10912 5220 11936
rect 4900 10848 4908 10912
rect 4972 10848 4988 10912
rect 5052 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5220 10912
rect 4900 9862 5220 10848
rect 4900 9824 4942 9862
rect 5178 9824 5220 9862
rect 4900 9760 4908 9824
rect 5212 9760 5220 9824
rect 4900 9626 4942 9760
rect 5178 9626 5220 9760
rect 4900 8736 5220 9626
rect 4900 8672 4908 8736
rect 4972 8672 4988 8736
rect 5052 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5220 8736
rect 4900 7648 5220 8672
rect 4900 7584 4908 7648
rect 4972 7584 4988 7648
rect 5052 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5220 7648
rect 4900 6560 5220 7584
rect 4900 6496 4908 6560
rect 4972 6496 4988 6560
rect 5052 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5220 6560
rect 4900 6054 5220 6496
rect 4900 5818 4942 6054
rect 5178 5818 5220 6054
rect 4900 5472 5220 5818
rect 4900 5408 4908 5472
rect 4972 5408 4988 5472
rect 5052 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5220 5472
rect 4900 4384 5220 5408
rect 4900 4320 4908 4384
rect 4972 4320 4988 4384
rect 5052 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5220 4384
rect 4900 3296 5220 4320
rect 4900 3232 4908 3296
rect 4972 3232 4988 3296
rect 5052 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5220 3296
rect 4900 2208 5220 3232
rect 4900 2144 4908 2208
rect 4972 2144 4988 2208
rect 5052 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5220 2208
rect 4900 2128 5220 2144
rect 6878 13632 7198 13648
rect 6878 13568 6886 13632
rect 6950 13568 6966 13632
rect 7030 13568 7046 13632
rect 7110 13568 7126 13632
rect 7190 13568 7198 13632
rect 6878 12544 7198 13568
rect 6878 12480 6886 12544
rect 6950 12480 6966 12544
rect 7030 12480 7046 12544
rect 7110 12480 7126 12544
rect 7190 12480 7198 12544
rect 6878 11766 7198 12480
rect 6878 11530 6920 11766
rect 7156 11530 7198 11766
rect 6878 11456 7198 11530
rect 6878 11392 6886 11456
rect 6950 11392 6966 11456
rect 7030 11392 7046 11456
rect 7110 11392 7126 11456
rect 7190 11392 7198 11456
rect 6878 10368 7198 11392
rect 6878 10304 6886 10368
rect 6950 10304 6966 10368
rect 7030 10304 7046 10368
rect 7110 10304 7126 10368
rect 7190 10304 7198 10368
rect 6878 9280 7198 10304
rect 6878 9216 6886 9280
rect 6950 9216 6966 9280
rect 7030 9216 7046 9280
rect 7110 9216 7126 9280
rect 7190 9216 7198 9280
rect 6878 8192 7198 9216
rect 6878 8128 6886 8192
rect 6950 8128 6966 8192
rect 7030 8128 7046 8192
rect 7110 8128 7126 8192
rect 7190 8128 7198 8192
rect 6878 7958 7198 8128
rect 6878 7722 6920 7958
rect 7156 7722 7198 7958
rect 6878 7104 7198 7722
rect 8856 13088 9176 13648
rect 8856 13024 8864 13088
rect 8928 13024 8944 13088
rect 9008 13024 9024 13088
rect 9088 13024 9104 13088
rect 9168 13024 9176 13088
rect 8856 12000 9176 13024
rect 8856 11936 8864 12000
rect 8928 11936 8944 12000
rect 9008 11936 9024 12000
rect 9088 11936 9104 12000
rect 9168 11936 9176 12000
rect 8856 10912 9176 11936
rect 8856 10848 8864 10912
rect 8928 10848 8944 10912
rect 9008 10848 9024 10912
rect 9088 10848 9104 10912
rect 9168 10848 9176 10912
rect 8856 9862 9176 10848
rect 8856 9824 8898 9862
rect 9134 9824 9176 9862
rect 8856 9760 8864 9824
rect 9168 9760 9176 9824
rect 8856 9626 8898 9760
rect 9134 9626 9176 9760
rect 8856 8736 9176 9626
rect 8856 8672 8864 8736
rect 8928 8672 8944 8736
rect 9008 8672 9024 8736
rect 9088 8672 9104 8736
rect 9168 8672 9176 8736
rect 8856 7648 9176 8672
rect 8856 7584 8864 7648
rect 8928 7584 8944 7648
rect 9008 7584 9024 7648
rect 9088 7584 9104 7648
rect 9168 7584 9176 7648
rect 7603 7172 7669 7173
rect 7603 7108 7604 7172
rect 7668 7108 7669 7172
rect 7603 7107 7669 7108
rect 6878 7040 6886 7104
rect 6950 7040 6966 7104
rect 7030 7040 7046 7104
rect 7110 7040 7126 7104
rect 7190 7040 7198 7104
rect 6878 6016 7198 7040
rect 6878 5952 6886 6016
rect 6950 5952 6966 6016
rect 7030 5952 7046 6016
rect 7110 5952 7126 6016
rect 7190 5952 7198 6016
rect 6878 4928 7198 5952
rect 7606 5677 7666 7107
rect 8856 6560 9176 7584
rect 8856 6496 8864 6560
rect 8928 6496 8944 6560
rect 9008 6496 9024 6560
rect 9088 6496 9104 6560
rect 9168 6496 9176 6560
rect 8856 6054 9176 6496
rect 10834 13632 11154 13648
rect 10834 13568 10842 13632
rect 10906 13568 10922 13632
rect 10986 13568 11002 13632
rect 11066 13568 11082 13632
rect 11146 13568 11154 13632
rect 10834 12544 11154 13568
rect 10834 12480 10842 12544
rect 10906 12480 10922 12544
rect 10986 12480 11002 12544
rect 11066 12480 11082 12544
rect 11146 12480 11154 12544
rect 10834 11766 11154 12480
rect 10834 11530 10876 11766
rect 11112 11530 11154 11766
rect 10834 11456 11154 11530
rect 10834 11392 10842 11456
rect 10906 11392 10922 11456
rect 10986 11392 11002 11456
rect 11066 11392 11082 11456
rect 11146 11392 11154 11456
rect 10834 10368 11154 11392
rect 10834 10304 10842 10368
rect 10906 10304 10922 10368
rect 10986 10304 11002 10368
rect 11066 10304 11082 10368
rect 11146 10304 11154 10368
rect 10834 9280 11154 10304
rect 10834 9216 10842 9280
rect 10906 9216 10922 9280
rect 10986 9216 11002 9280
rect 11066 9216 11082 9280
rect 11146 9216 11154 9280
rect 10834 8192 11154 9216
rect 10834 8128 10842 8192
rect 10906 8128 10922 8192
rect 10986 8128 11002 8192
rect 11066 8128 11082 8192
rect 11146 8128 11154 8192
rect 10834 7958 11154 8128
rect 10834 7722 10876 7958
rect 11112 7722 11154 7958
rect 10834 7104 11154 7722
rect 10834 7040 10842 7104
rect 10906 7040 10922 7104
rect 10986 7040 11002 7104
rect 11066 7040 11082 7104
rect 11146 7040 11154 7104
rect 9995 6492 10061 6493
rect 9995 6428 9996 6492
rect 10060 6428 10061 6492
rect 9995 6427 10061 6428
rect 8856 5818 8898 6054
rect 9134 5818 9176 6054
rect 7603 5676 7669 5677
rect 7603 5612 7604 5676
rect 7668 5612 7669 5676
rect 7603 5611 7669 5612
rect 6878 4864 6886 4928
rect 6950 4864 6966 4928
rect 7030 4864 7046 4928
rect 7110 4864 7126 4928
rect 7190 4864 7198 4928
rect 6878 4150 7198 4864
rect 6878 3914 6920 4150
rect 7156 3914 7198 4150
rect 6878 3840 7198 3914
rect 6878 3776 6886 3840
rect 6950 3776 6966 3840
rect 7030 3776 7046 3840
rect 7110 3776 7126 3840
rect 7190 3776 7198 3840
rect 6878 2752 7198 3776
rect 6878 2688 6886 2752
rect 6950 2688 6966 2752
rect 7030 2688 7046 2752
rect 7110 2688 7126 2752
rect 7190 2688 7198 2752
rect 6878 2128 7198 2688
rect 8856 5472 9176 5818
rect 8856 5408 8864 5472
rect 8928 5408 8944 5472
rect 9008 5408 9024 5472
rect 9088 5408 9104 5472
rect 9168 5408 9176 5472
rect 8856 4384 9176 5408
rect 8856 4320 8864 4384
rect 8928 4320 8944 4384
rect 9008 4320 9024 4384
rect 9088 4320 9104 4384
rect 9168 4320 9176 4384
rect 8856 3296 9176 4320
rect 9998 4045 10058 6427
rect 10834 6016 11154 7040
rect 10834 5952 10842 6016
rect 10906 5952 10922 6016
rect 10986 5952 11002 6016
rect 11066 5952 11082 6016
rect 11146 5952 11154 6016
rect 10834 4928 11154 5952
rect 10834 4864 10842 4928
rect 10906 4864 10922 4928
rect 10986 4864 11002 4928
rect 11066 4864 11082 4928
rect 11146 4864 11154 4928
rect 10834 4150 11154 4864
rect 9995 4044 10061 4045
rect 9995 3980 9996 4044
rect 10060 3980 10061 4044
rect 9995 3979 10061 3980
rect 8856 3232 8864 3296
rect 8928 3232 8944 3296
rect 9008 3232 9024 3296
rect 9088 3232 9104 3296
rect 9168 3232 9176 3296
rect 8856 2208 9176 3232
rect 8856 2144 8864 2208
rect 8928 2144 8944 2208
rect 9008 2144 9024 2208
rect 9088 2144 9104 2208
rect 9168 2144 9176 2208
rect 8856 2128 9176 2144
rect 10834 3914 10876 4150
rect 11112 3914 11154 4150
rect 10834 3840 11154 3914
rect 10834 3776 10842 3840
rect 10906 3776 10922 3840
rect 10986 3776 11002 3840
rect 11066 3776 11082 3840
rect 11146 3776 11154 3840
rect 10834 2752 11154 3776
rect 10834 2688 10842 2752
rect 10906 2688 10922 2752
rect 10986 2688 11002 2752
rect 11066 2688 11082 2752
rect 11146 2688 11154 2752
rect 10834 2128 11154 2688
<< via4 >>
rect 2964 11530 3200 11766
rect 2964 7722 3200 7958
rect 2964 3914 3200 4150
rect 4942 9824 5178 9862
rect 4942 9760 4972 9824
rect 4972 9760 4988 9824
rect 4988 9760 5052 9824
rect 5052 9760 5068 9824
rect 5068 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5178 9824
rect 4942 9626 5178 9760
rect 4942 5818 5178 6054
rect 6920 11530 7156 11766
rect 6920 7722 7156 7958
rect 8898 9824 9134 9862
rect 8898 9760 8928 9824
rect 8928 9760 8944 9824
rect 8944 9760 9008 9824
rect 9008 9760 9024 9824
rect 9024 9760 9088 9824
rect 9088 9760 9104 9824
rect 9104 9760 9134 9824
rect 8898 9626 9134 9760
rect 10876 11530 11112 11766
rect 10876 7722 11112 7958
rect 8898 5818 9134 6054
rect 6920 3914 7156 4150
rect 10876 3914 11112 4150
<< metal5 >>
rect 1104 11766 12972 11808
rect 1104 11530 2964 11766
rect 3200 11530 6920 11766
rect 7156 11530 10876 11766
rect 11112 11530 12972 11766
rect 1104 11488 12972 11530
rect 1104 9862 12972 9904
rect 1104 9626 4942 9862
rect 5178 9626 8898 9862
rect 9134 9626 12972 9862
rect 1104 9584 12972 9626
rect 1104 7958 12972 8000
rect 1104 7722 2964 7958
rect 3200 7722 6920 7958
rect 7156 7722 10876 7958
rect 11112 7722 12972 7958
rect 1104 7680 12972 7722
rect 1104 6054 12972 6096
rect 1104 5818 4942 6054
rect 5178 5818 8898 6054
rect 9134 5818 12972 6054
rect 1104 5776 12972 5818
rect 1104 4150 12972 4192
rect 1104 3914 2964 4150
rect 3200 3914 6920 4150
rect 7156 3914 10876 4150
rect 11112 3914 12972 4150
rect 1104 3872 12972 3914
use sky130_fd_sc_hd__decap_6  FILLER_0_11
timestamp 1630053115
transform 1 0 2116 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1630053115
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_6
timestamp 1630053115
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1630053115
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1630053115
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1630053115
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output27
timestamp 1630053115
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21
timestamp 1630053115
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_18
timestamp 1630053115
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output28
timestamp 1630053115
transform -1 0 3036 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1630053115
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1630053115
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34
timestamp 1630053115
transform 1 0 4232 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_30
timestamp 1630053115
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1630053115
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1630053115
transform 1 0 3956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42
timestamp 1630053115
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49
timestamp 1630053115
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_42
timestamp 1630053115
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output31
timestamp 1630053115
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1630053115
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1630053115
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62
timestamp 1630053115
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1630053115
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1630053115
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1630053115
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1630053115
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1630053115
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1630053115
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1630053115
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1630053115
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1630053115
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1630053115
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output36
timestamp 1630053115
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1630053115
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1630053115
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_86
timestamp 1630053115
transform 1 0 9016 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1630053115
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _112_
timestamp 1630053115
transform -1 0 9016 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1630053115
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1630053115
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_90
timestamp 1630053115
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1630053115
transform 1 0 9568 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__dlxtp_1  _123_
timestamp 1630053115
transform -1 0 10764 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1630053115
transform -1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1630053115
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1630053115
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1630053115
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1630053115
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1630053115
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1630053115
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1630053115
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1630053115
transform 1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1630053115
transform -1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_117
timestamp 1630053115
transform 1 0 11868 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1630053115
transform 1 0 12604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_117
timestamp 1630053115
transform 1 0 11868 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_122
timestamp 1630053115
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1630053115
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1630053115
transform -1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output30
timestamp 1630053115
transform 1 0 11960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_6
timestamp 1630053115
transform 1 0 1656 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1630053115
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1630053115
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_18
timestamp 1630053115
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1630053115
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1630053115
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1630053115
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1630053115
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_53
timestamp 1630053115
transform 1 0 5980 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2oi_1  _109_
timestamp 1630053115
transform -1 0 7360 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1630053115
transform 1 0 7360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1630053115
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_85
timestamp 1630053115
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1630053115
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 1630053115
transform 1 0 9476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1630053115
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _115_
timestamp 1630053115
transform -1 0 10212 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_2_106
timestamp 1630053115
transform 1 0 10856 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _064_
timestamp 1630053115
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1630053115
transform -1 0 12328 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1630053115
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1630053115
transform -1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_11
timestamp 1630053115
transform 1 0 2116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1630053115
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1630053115
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output29
timestamp 1630053115
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_23
timestamp 1630053115
transform 1 0 3220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_29
timestamp 1630053115
transform 1 0 3772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_33
timestamp 1630053115
transform 1 0 4140 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _068_
timestamp 1630053115
transform -1 0 4140 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1630053115
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1630053115
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1630053115
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1630053115
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_69
timestamp 1630053115
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_77
timestamp 1630053115
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_88
timestamp 1630053115
transform 1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _101_
timestamp 1630053115
transform -1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_99
timestamp 1630053115
transform 1 0 10212 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1630053115
transform -1 0 10212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1630053115
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1630053115
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1630053115
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _087_
timestamp 1630053115
transform 1 0 11684 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _100_
timestamp 1630053115
transform 1 0 10580 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_3_120
timestamp 1630053115
transform 1 0 12144 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1630053115
transform -1 0 12972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1630053115
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1630053115
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1630053115
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _106_
timestamp 1630053115
transform 1 0 2024 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_18
timestamp 1630053115
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1630053115
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_36
timestamp 1630053115
transform 1 0 4416 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1630053115
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _084_
timestamp 1630053115
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlxtp_1  _124_
timestamp 1630053115
transform -1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1630053115
transform 1 0 6072 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1630053115
transform 1 0 7176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1630053115
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1630053115
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1630053115
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1630053115
transform -1 0 9568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_92
timestamp 1630053115
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_104
timestamp 1630053115
transform 1 0 10672 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _072_
timestamp 1630053115
transform -1 0 11868 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_4_117
timestamp 1630053115
transform 1 0 11868 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1630053115
transform 1 0 12604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1630053115
transform -1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1630053115
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1630053115
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1630053115
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _095_
timestamp 1630053115
transform 1 0 3220 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_5_30
timestamp 1630053115
transform 1 0 3864 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_42
timestamp 1630053115
transform 1 0 4968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1630053115
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1630053115
transform -1 0 5336 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1630053115
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_60
timestamp 1630053115
transform 1 0 6624 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1630053115
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _062_
timestamp 1630053115
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_72
timestamp 1630053115
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1630053115
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_96
timestamp 1630053115
transform 1 0 9936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1630053115
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1630053115
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1630053115
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _081_
timestamp 1630053115
transform 1 0 11684 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_122
timestamp 1630053115
transform 1 0 12328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1630053115
transform -1 0 12972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1630053115
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_6
timestamp 1630053115
transform 1 0 1656 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1630053115
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1630053115
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1630053115
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1630053115
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1630053115
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_23
timestamp 1630053115
transform 1 0 3220 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_1  _097_
timestamp 1630053115
transform 1 0 2576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1630053115
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1630053115
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1630053115
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1630053115
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _085_
timestamp 1630053115
transform 1 0 4324 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _093_
timestamp 1630053115
transform -1 0 5060 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1630053115
transform 1 0 5060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1630053115
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _117_
timestamp 1630053115
transform -1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_59
timestamp 1630053115
transform 1 0 6532 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1630053115
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1630053115
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1630053115
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _105_
timestamp 1630053115
transform -1 0 7544 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_6_70
timestamp 1630053115
transform 1 0 7544 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1630053115
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_73
timestamp 1630053115
transform 1 0 7820 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _066_
timestamp 1630053115
transform -1 0 7820 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1630053115
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_85
timestamp 1630053115
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp 1630053115
transform 1 0 8924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_89
timestamp 1630053115
transform 1 0 9292 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1630053115
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 1630053115
transform -1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1630053115
transform 1 0 9660 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__dlxtp_1  _120_
timestamp 1630053115
transform -1 0 10764 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _126_
timestamp 1630053115
transform -1 0 10948 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_107
timestamp 1630053115
transform 1 0 10948 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_115
timestamp 1630053115
transform 1 0 11684 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1630053115
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1630053115
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1630053115
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _102_
timestamp 1630053115
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_121
timestamp 1630053115
transform 1 0 12236 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_125
timestamp 1630053115
transform 1 0 12604 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_121
timestamp 1630053115
transform 1 0 12236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_125
timestamp 1630053115
transform 1 0 12604 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1630053115
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1630053115
transform -1 0 12972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 1630053115
transform -1 0 12236 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1630053115
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1630053115
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtp_1  _118_
timestamp 1630053115
transform -1 0 2576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_16
timestamp 1630053115
transform 1 0 2576 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1630053115
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1630053115
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1630053115
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1630053115
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1630053115
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _075_
timestamp 1630053115
transform -1 0 6808 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_8_73
timestamp 1630053115
transform 1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _060_
timestamp 1630053115
transform 1 0 7176 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_8_81
timestamp 1630053115
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1630053115
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1630053115
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1630053115
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 1630053115
transform 1 0 11132 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_117
timestamp 1630053115
transform 1 0 11868 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1630053115
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1630053115
transform -1 0 12972 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output39
timestamp 1630053115
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1630053115
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1630053115
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp 1630053115
transform -1 0 2300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1630053115
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_13
timestamp 1630053115
transform 1 0 2300 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlxtp_1  _122_
timestamp 1630053115
transform 1 0 2852 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_31
timestamp 1630053115
transform 1 0 3956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_43
timestamp 1630053115
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1630053115
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1630053115
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1630053115
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_65
timestamp 1630053115
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_75
timestamp 1630053115
transform 1 0 8004 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _108_
timestamp 1630053115
transform -1 0 8004 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1630053115
transform 1 0 8648 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _071_
timestamp 1630053115
transform -1 0 8648 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1630053115
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1630053115
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1630053115
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1630053115
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_125
timestamp 1630053115
transform 1 0 12604 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1630053115
transform -1 0 12972 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1630053115
transform 1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1630053115
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2oi_1  _110_
timestamp 1630053115
transform 1 0 2116 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  output37
timestamp 1630053115
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_18
timestamp 1630053115
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1630053115
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1630053115
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1630053115
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1630053115
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1630053115
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1630053115
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1630053115
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1630053115
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1630053115
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1630053115
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1630053115
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_109
timestamp 1630053115
transform 1 0 11132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1630053115
transform -1 0 12328 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_10_122
timestamp 1630053115
transform 1 0 12328 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1630053115
transform -1 0 12972 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1630053115
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1630053115
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1630053115
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1630053115
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1630053115
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1630053115
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1630053115
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1630053115
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1630053115
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_69
timestamp 1630053115
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_73
timestamp 1630053115
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlxtp_1  _128_
timestamp 1630053115
transform -1 0 9016 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_86
timestamp 1630053115
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_97
timestamp 1630053115
transform 1 0 10028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__a22o_1  _078_
timestamp 1630053115
transform -1 0 10028 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1630053115
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1630053115
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1630053115
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_125
timestamp 1630053115
transform 1 0 12604 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1630053115
transform -1 0 12972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1630053115
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1630053115
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1630053115
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtp_1  _127_
timestamp 1630053115
transform 1 0 1840 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_20
timestamp 1630053115
transform 1 0 2944 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1630053115
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1630053115
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__dlxtp_1  _121_
timestamp 1630053115
transform 1 0 4048 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_44
timestamp 1630053115
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _096_
timestamp 1630053115
transform 1 0 5520 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_55
timestamp 1630053115
transform 1 0 6164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_67
timestamp 1630053115
transform 1 0 7268 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1630053115
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1630053115
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1630053115
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1630053115
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_101
timestamp 1630053115
transform 1 0 10396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1630053115
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _063_
timestamp 1630053115
transform -1 0 10396 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_113
timestamp 1630053115
transform 1 0 11500 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_125
timestamp 1630053115
transform 1 0 12604 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1630053115
transform -1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1630053115
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_11
timestamp 1630053115
transform 1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1630053115
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1630053115
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1630053115
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1630053115
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1630053115
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_18
timestamp 1630053115
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1630053115
transform -1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1630053115
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1630053115
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_29
timestamp 1630053115
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_38
timestamp 1630053115
transform 1 0 4600 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1630053115
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _067_
timestamp 1630053115
transform -1 0 4600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1630053115
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1630053115
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_50
timestamp 1630053115
transform 1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1630053115
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1630053115
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_63
timestamp 1630053115
transform 1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1630053115
transform 1 0 6808 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1630053115
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1630053115
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_69
timestamp 1630053115
transform 1 0 7452 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_74
timestamp 1630053115
transform 1 0 7912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlxtp_1  _116_
timestamp 1630053115
transform -1 0 8648 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1630053115
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1630053115
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1630053115
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__a22o_1  _069_
timestamp 1630053115
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlxtp_1  _119_
timestamp 1630053115
transform 1 0 9016 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1630053115
transform 1 0 10120 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1630053115
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_99
timestamp 1630053115
transform 1 0 10212 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _061_
timestamp 1630053115
transform 1 0 9936 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1630053115
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1630053115
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_110
timestamp 1630053115
transform 1 0 11224 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1630053115
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1630053115
transform 1 0 10948 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_125
timestamp 1630053115
transform 1 0 12604 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_118
timestamp 1630053115
transform 1 0 11960 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_122
timestamp 1630053115
transform 1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1630053115
transform -1 0 12972 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1630053115
transform -1 0 12972 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1630053115
transform -1 0 12328 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1630053115
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1630053115
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1630053115
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1630053115
transform 1 0 3588 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1630053115
transform 1 0 4416 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _103_
timestamp 1630053115
transform 1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1630053115
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _088_
timestamp 1630053115
transform -1 0 5428 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1630053115
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1630053115
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1630053115
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1630053115
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1630053115
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1630053115
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1630053115
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1630053115
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1630053115
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1630053115
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_125
timestamp 1630053115
transform 1 0 12604 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1630053115
transform -1 0 12972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1630053115
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1630053115
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1630053115
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1630053115
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1630053115
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1630053115
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1630053115
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 1630053115
transform -1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1630053115
transform 1 0 4876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp 1630053115
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_1  _092_
timestamp 1630053115
transform -1 0 6440 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_16_58
timestamp 1630053115
transform 1 0 6440 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_70
timestamp 1630053115
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1630053115
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1630053115
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1630053115
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_97
timestamp 1630053115
transform 1 0 10028 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_105
timestamp 1630053115
transform 1 0 10764 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_115
timestamp 1630053115
transform 1 0 11684 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _107_
timestamp 1630053115
transform -1 0 11684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1630053115
transform 1 0 12328 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1630053115
transform -1 0 12972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1630053115
transform -1 0 12328 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1630053115
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1630053115
transform 1 0 1380 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1630053115
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1630053115
transform 1 0 2668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1630053115
transform 1 0 3404 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2oi_1  _114_
timestamp 1630053115
transform 1 0 2760 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1630053115
transform 1 0 4508 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_49
timestamp 1630053115
transform 1 0 5612 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1630053115
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_64
timestamp 1630053115
transform 1 0 6992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1630053115
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _094_
timestamp 1630053115
transform 1 0 6348 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_17_76
timestamp 1630053115
transform 1 0 8096 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_88
timestamp 1630053115
transform 1 0 9200 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1630053115
transform 1 0 10396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1630053115
transform 1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1630053115
transform -1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1630053115
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1630053115
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1630053115
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _082_
timestamp 1630053115
transform 1 0 10764 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _098_
timestamp 1630053115
transform -1 0 12328 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_122
timestamp 1630053115
transform 1 0 12328 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1630053115
transform -1 0 12972 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1630053115
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtp_1  _125_
timestamp 1630053115
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1630053115
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1630053115
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_36
timestamp 1630053115
transform 1 0 4416 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1630053115
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _111_
timestamp 1630053115
transform 1 0 3772 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_18_48
timestamp 1630053115
transform 1 0 5520 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_60
timestamp 1630053115
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_72
timestamp 1630053115
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_85
timestamp 1630053115
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1630053115
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_96
timestamp 1630053115
transform 1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1630053115
transform -1 0 9936 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1630053115
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1630053115
transform -1 0 12328 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  output33
timestamp 1630053115
transform 1 0 10672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_122
timestamp 1630053115
transform 1 0 12328 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1630053115
transform -1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_11
timestamp 1630053115
transform 1 0 2116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1630053115
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_11
timestamp 1630053115
transform 1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1630053115
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1630053115
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1630053115
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output32
timestamp 1630053115
transform -1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output38
timestamp 1630053115
transform -1 0 2116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1630053115
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _080_
timestamp 1630053115
transform -1 0 3496 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1630053115
transform 1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_26
timestamp 1630053115
transform 1 0 3496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1630053115
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1630053115
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1630053115
transform 1 0 4048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1630053115
transform 1 0 4416 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1630053115
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2oi_1  _113_
timestamp 1630053115
transform -1 0 4508 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1630053115
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1630053115
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1630053115
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 1630053115
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_47
timestamp 1630053115
transform 1 0 5428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1630053115
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1630053115
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_57
timestamp 1630053115
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_61
timestamp 1630053115
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_55
timestamp 1630053115
transform 1 0 6164 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_57
timestamp 1630053115
transform 1 0 6348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1630053115
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1630053115
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__a31oi_2  _091_
timestamp 1630053115
transform 1 0 6808 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  output34
timestamp 1630053115
transform -1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_72
timestamp 1630053115
transform 1 0 7728 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1630053115
transform 1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_73
timestamp 1630053115
transform 1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1630053115
transform -1 0 8464 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output35
timestamp 1630053115
transform -1 0 7820 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_84
timestamp 1630053115
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1630053115
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1630053115
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1630053115
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _089_
timestamp 1630053115
transform 1 0 9292 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _099_
timestamp 1630053115
transform -1 0 9660 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1630053115
transform 1 0 10396 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_93
timestamp 1630053115
transform 1 0 9660 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1630053115
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1630053115
transform -1 0 11040 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input25
timestamp 1630053115
transform -1 0 11040 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1630053115
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_108
timestamp 1630053115
transform 1 0 11040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1630053115
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1630053115
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__o2bb2a_1  _086_
timestamp 1630053115
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _090_
timestamp 1630053115
transform 1 0 11500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_121
timestamp 1630053115
transform 1 0 12236 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_125
timestamp 1630053115
transform 1 0 12604 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_121
timestamp 1630053115
transform 1 0 12236 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_125
timestamp 1630053115
transform 1 0 12604 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1630053115
transform -1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1630053115
transform -1 0 12972 0 1 13056
box -38 -48 314 592
<< labels >>
rlabel metal2 s 9034 0 9090 800 4 A[0]
port 1 nsew
rlabel metal2 s 6458 0 6514 800 4 A[10]
port 2 nsew
rlabel metal2 s 9586 15506 9642 16306 4 A[11]
port 3 nsew
rlabel metal3 s 13362 7624 14162 7744 4 A[1]
port 4 nsew
rlabel metal3 s 0 5720 800 5840 4 A[2]
port 5 nsew
rlabel metal2 s 8298 15506 8354 16306 4 A[3]
port 6 nsew
rlabel metal2 s 12898 0 12954 800 4 A[4]
port 7 nsew
rlabel metal2 s 3146 15506 3202 16306 4 A[5]
port 8 nsew
rlabel metal3 s 13362 11432 14162 11552 4 A[6]
port 9 nsew
rlabel metal2 s 11610 0 11666 800 4 A[7]
port 10 nsew
rlabel metal2 s 13450 15506 13506 16306 4 A[8]
port 11 nsew
rlabel metal3 s 13362 13336 14162 13456 4 A[9]
port 12 nsew
rlabel metal2 s 4434 15506 4490 16306 4 B[0]
port 13 nsew
rlabel metal3 s 0 15240 800 15360 4 B[10]
port 14 nsew
rlabel metal3 s 13362 1912 14162 2032 4 B[11]
port 15 nsew
rlabel metal3 s 0 9528 800 9648 4 B[1]
port 16 nsew
rlabel metal3 s 13362 9528 14162 9648 4 B[2]
port 17 nsew
rlabel metal3 s 0 11432 800 11552 4 B[3]
port 18 nsew
rlabel metal2 s 18 0 74 800 4 B[4]
port 19 nsew
rlabel metal2 s 10874 15506 10930 16306 4 B[5]
port 20 nsew
rlabel metal3 s 0 1912 800 2032 4 B[6]
port 21 nsew
rlabel metal2 s 3882 0 3938 800 4 B[7]
port 22 nsew
rlabel metal2 s 1858 15506 1914 16306 4 B[8]
port 23 nsew
rlabel metal2 s 10322 0 10378 800 4 B[9]
port 24 nsew
rlabel metal2 s 12162 15506 12218 16306 4 CE
port 25 nsew
rlabel metal3 s 13362 8 14162 128 4 Cin
port 26 nsew
rlabel metal2 s 1306 0 1362 800 4 Cout
port 27 nsew
rlabel metal2 s 2594 0 2650 800 4 S[0]
port 28 nsew
rlabel metal3 s 0 3816 800 3936 4 S[10]
port 29 nsew
rlabel metal3 s 13362 3816 14162 3936 4 S[11]
port 30 nsew
rlabel metal2 s 5170 0 5226 800 4 S[1]
port 31 nsew
rlabel metal3 s 0 13336 800 13456 4 S[2]
port 32 nsew
rlabel metal3 s 13362 15240 14162 15360 4 S[3]
port 33 nsew
rlabel metal2 s 5722 15506 5778 16306 4 S[4]
port 34 nsew
rlabel metal2 s 7010 15506 7066 16306 4 S[5]
port 35 nsew
rlabel metal2 s 7746 0 7802 800 4 S[6]
port 36 nsew
rlabel metal3 s 0 7624 800 7744 4 S[7]
port 37 nsew
rlabel metal2 s 570 15506 626 16306 4 S[8]
port 38 nsew
rlabel metal3 s 13362 5720 14162 5840 4 S[9]
port 39 nsew
rlabel metal5 s 1104 5776 12972 6096 4 VGND
port 40 nsew
rlabel metal5 s 1104 3872 12972 4192 4 VPWR
port 41 nsew
<< properties >>
string FIXED_BBOX 0 0 14162 16306
<< end >>
